
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"d8",x"df",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"d8",x"df",x"c2"),
    14 => (x"48",x"d8",x"cd",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"d5",x"dc"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d6",x"02",x"99"),
    50 => (x"c3",x"48",x"d4",x"ff"),
    51 => (x"52",x"68",x"78",x"ff"),
    52 => (x"48",x"49",x"66",x"c4"),
    53 => (x"a6",x"c8",x"88",x"c1"),
    54 => (x"05",x"99",x"71",x"58"),
    55 => (x"4f",x"26",x"87",x"ea"),
    56 => (x"ff",x"1e",x"73",x"1e"),
    57 => (x"ff",x"c3",x"4b",x"d4"),
    58 => (x"c3",x"4a",x"6b",x"7b"),
    59 => (x"49",x"6b",x"7b",x"ff"),
    60 => (x"b1",x"72",x"32",x"c8"),
    61 => (x"6b",x"7b",x"ff",x"c3"),
    62 => (x"71",x"31",x"c8",x"4a"),
    63 => (x"7b",x"ff",x"c3",x"b2"),
    64 => (x"32",x"c8",x"49",x"6b"),
    65 => (x"48",x"71",x"b1",x"72"),
    66 => (x"4d",x"26",x"87",x"c4"),
    67 => (x"4b",x"26",x"4c",x"26"),
    68 => (x"5e",x"0e",x"4f",x"26"),
    69 => (x"0e",x"5d",x"5c",x"5b"),
    70 => (x"d4",x"ff",x"4a",x"71"),
    71 => (x"c3",x"48",x"72",x"4c"),
    72 => (x"7c",x"70",x"98",x"ff"),
    73 => (x"bf",x"d8",x"cd",x"c2"),
    74 => (x"d0",x"87",x"c8",x"05"),
    75 => (x"30",x"c9",x"48",x"66"),
    76 => (x"d0",x"58",x"a6",x"d4"),
    77 => (x"29",x"d8",x"49",x"66"),
    78 => (x"ff",x"c3",x"48",x"71"),
    79 => (x"d0",x"7c",x"70",x"98"),
    80 => (x"29",x"d0",x"49",x"66"),
    81 => (x"71",x"99",x"ff",x"c3"),
    82 => (x"49",x"66",x"d0",x"7c"),
    83 => (x"ff",x"c3",x"29",x"c8"),
    84 => (x"d0",x"7c",x"71",x"99"),
    85 => (x"ff",x"c3",x"49",x"66"),
    86 => (x"72",x"7c",x"71",x"99"),
    87 => (x"71",x"29",x"d0",x"49"),
    88 => (x"98",x"ff",x"c3",x"48"),
    89 => (x"4b",x"6c",x"7c",x"70"),
    90 => (x"4d",x"ff",x"f0",x"c9"),
    91 => (x"05",x"ab",x"ff",x"c3"),
    92 => (x"ff",x"c3",x"87",x"d0"),
    93 => (x"c1",x"4b",x"6c",x"7c"),
    94 => (x"87",x"c6",x"02",x"8d"),
    95 => (x"02",x"ab",x"ff",x"c3"),
    96 => (x"48",x"73",x"87",x"f0"),
    97 => (x"1e",x"87",x"c3",x"fe"),
    98 => (x"d4",x"ff",x"49",x"c0"),
    99 => (x"78",x"ff",x"c3",x"48"),
   100 => (x"c8",x"c3",x"81",x"c1"),
   101 => (x"f1",x"04",x"a9",x"b7"),
   102 => (x"1e",x"4f",x"26",x"87"),
   103 => (x"87",x"e7",x"1e",x"73"),
   104 => (x"4b",x"df",x"f8",x"c4"),
   105 => (x"ff",x"c0",x"1e",x"c0"),
   106 => (x"49",x"f7",x"c1",x"f0"),
   107 => (x"c4",x"87",x"e3",x"fd"),
   108 => (x"05",x"a8",x"c1",x"86"),
   109 => (x"ff",x"87",x"ea",x"c0"),
   110 => (x"ff",x"c3",x"48",x"d4"),
   111 => (x"c0",x"c0",x"c1",x"78"),
   112 => (x"1e",x"c0",x"c0",x"c0"),
   113 => (x"c1",x"f0",x"e1",x"c0"),
   114 => (x"c5",x"fd",x"49",x"e9"),
   115 => (x"70",x"86",x"c4",x"87"),
   116 => (x"87",x"ca",x"05",x"98"),
   117 => (x"c3",x"48",x"d4",x"ff"),
   118 => (x"48",x"c1",x"78",x"ff"),
   119 => (x"e6",x"fe",x"87",x"cb"),
   120 => (x"05",x"8b",x"c1",x"87"),
   121 => (x"c0",x"87",x"fd",x"fe"),
   122 => (x"87",x"e2",x"fc",x"48"),
   123 => (x"ff",x"1e",x"73",x"1e"),
   124 => (x"ff",x"c3",x"48",x"d4"),
   125 => (x"c0",x"4b",x"d3",x"78"),
   126 => (x"f0",x"ff",x"c0",x"1e"),
   127 => (x"fc",x"49",x"c1",x"c1"),
   128 => (x"86",x"c4",x"87",x"d0"),
   129 => (x"ca",x"05",x"98",x"70"),
   130 => (x"48",x"d4",x"ff",x"87"),
   131 => (x"c1",x"78",x"ff",x"c3"),
   132 => (x"fd",x"87",x"cb",x"48"),
   133 => (x"8b",x"c1",x"87",x"f1"),
   134 => (x"87",x"db",x"ff",x"05"),
   135 => (x"ed",x"fb",x"48",x"c0"),
   136 => (x"5b",x"5e",x"0e",x"87"),
   137 => (x"d4",x"ff",x"0e",x"5c"),
   138 => (x"87",x"db",x"fd",x"4c"),
   139 => (x"c0",x"1e",x"ea",x"c6"),
   140 => (x"c8",x"c1",x"f0",x"e1"),
   141 => (x"87",x"da",x"fb",x"49"),
   142 => (x"a8",x"c1",x"86",x"c4"),
   143 => (x"fe",x"87",x"c8",x"02"),
   144 => (x"48",x"c0",x"87",x"ea"),
   145 => (x"fa",x"87",x"e2",x"c1"),
   146 => (x"49",x"70",x"87",x"d6"),
   147 => (x"99",x"ff",x"ff",x"cf"),
   148 => (x"02",x"a9",x"ea",x"c6"),
   149 => (x"d3",x"fe",x"87",x"c8"),
   150 => (x"c1",x"48",x"c0",x"87"),
   151 => (x"ff",x"c3",x"87",x"cb"),
   152 => (x"4b",x"f1",x"c0",x"7c"),
   153 => (x"70",x"87",x"f4",x"fc"),
   154 => (x"eb",x"c0",x"02",x"98"),
   155 => (x"c0",x"1e",x"c0",x"87"),
   156 => (x"fa",x"c1",x"f0",x"ff"),
   157 => (x"87",x"da",x"fa",x"49"),
   158 => (x"98",x"70",x"86",x"c4"),
   159 => (x"c3",x"87",x"d9",x"05"),
   160 => (x"49",x"6c",x"7c",x"ff"),
   161 => (x"7c",x"7c",x"ff",x"c3"),
   162 => (x"c0",x"c1",x"7c",x"7c"),
   163 => (x"87",x"c4",x"02",x"99"),
   164 => (x"87",x"d5",x"48",x"c1"),
   165 => (x"87",x"d1",x"48",x"c0"),
   166 => (x"c4",x"05",x"ab",x"c2"),
   167 => (x"c8",x"48",x"c0",x"87"),
   168 => (x"05",x"8b",x"c1",x"87"),
   169 => (x"c0",x"87",x"fd",x"fe"),
   170 => (x"87",x"e0",x"f9",x"48"),
   171 => (x"c2",x"1e",x"73",x"1e"),
   172 => (x"c1",x"48",x"d8",x"cd"),
   173 => (x"ff",x"4b",x"c7",x"78"),
   174 => (x"78",x"c2",x"48",x"d0"),
   175 => (x"ff",x"87",x"c8",x"fb"),
   176 => (x"78",x"c3",x"48",x"d0"),
   177 => (x"e5",x"c0",x"1e",x"c0"),
   178 => (x"49",x"c0",x"c1",x"d0"),
   179 => (x"c4",x"87",x"c3",x"f9"),
   180 => (x"05",x"a8",x"c1",x"86"),
   181 => (x"c2",x"4b",x"87",x"c1"),
   182 => (x"87",x"c5",x"05",x"ab"),
   183 => (x"f9",x"c0",x"48",x"c0"),
   184 => (x"05",x"8b",x"c1",x"87"),
   185 => (x"fc",x"87",x"d0",x"ff"),
   186 => (x"cd",x"c2",x"87",x"f7"),
   187 => (x"98",x"70",x"58",x"dc"),
   188 => (x"c1",x"87",x"cd",x"05"),
   189 => (x"f0",x"ff",x"c0",x"1e"),
   190 => (x"f8",x"49",x"d0",x"c1"),
   191 => (x"86",x"c4",x"87",x"d4"),
   192 => (x"c3",x"48",x"d4",x"ff"),
   193 => (x"fd",x"c2",x"78",x"ff"),
   194 => (x"e0",x"cd",x"c2",x"87"),
   195 => (x"48",x"d0",x"ff",x"58"),
   196 => (x"d4",x"ff",x"78",x"c2"),
   197 => (x"78",x"ff",x"c3",x"48"),
   198 => (x"f1",x"f7",x"48",x"c1"),
   199 => (x"5b",x"5e",x"0e",x"87"),
   200 => (x"71",x"0e",x"5d",x"5c"),
   201 => (x"c5",x"4c",x"c0",x"4b"),
   202 => (x"4a",x"df",x"cd",x"ee"),
   203 => (x"c3",x"48",x"d4",x"ff"),
   204 => (x"48",x"68",x"78",x"ff"),
   205 => (x"05",x"a8",x"fe",x"c3"),
   206 => (x"ff",x"87",x"fe",x"c0"),
   207 => (x"9b",x"73",x"4d",x"d4"),
   208 => (x"d0",x"87",x"cc",x"02"),
   209 => (x"49",x"73",x"1e",x"66"),
   210 => (x"c4",x"87",x"ec",x"f5"),
   211 => (x"ff",x"87",x"d6",x"86"),
   212 => (x"d1",x"c4",x"48",x"d0"),
   213 => (x"7d",x"ff",x"c3",x"78"),
   214 => (x"c1",x"48",x"66",x"d0"),
   215 => (x"58",x"a6",x"d4",x"88"),
   216 => (x"f0",x"05",x"98",x"70"),
   217 => (x"48",x"d4",x"ff",x"87"),
   218 => (x"78",x"78",x"ff",x"c3"),
   219 => (x"c5",x"05",x"9b",x"73"),
   220 => (x"48",x"d0",x"ff",x"87"),
   221 => (x"4a",x"c1",x"78",x"d0"),
   222 => (x"05",x"8a",x"c1",x"4c"),
   223 => (x"74",x"87",x"ed",x"fe"),
   224 => (x"87",x"c6",x"f6",x"48"),
   225 => (x"71",x"1e",x"73",x"1e"),
   226 => (x"ff",x"4b",x"c0",x"4a"),
   227 => (x"ff",x"c3",x"48",x"d4"),
   228 => (x"48",x"d0",x"ff",x"78"),
   229 => (x"ff",x"78",x"c3",x"c4"),
   230 => (x"ff",x"c3",x"48",x"d4"),
   231 => (x"c0",x"1e",x"72",x"78"),
   232 => (x"d1",x"c1",x"f0",x"ff"),
   233 => (x"87",x"ea",x"f5",x"49"),
   234 => (x"98",x"70",x"86",x"c4"),
   235 => (x"c8",x"87",x"d2",x"05"),
   236 => (x"66",x"cc",x"1e",x"c0"),
   237 => (x"87",x"e5",x"fd",x"49"),
   238 => (x"4b",x"70",x"86",x"c4"),
   239 => (x"c2",x"48",x"d0",x"ff"),
   240 => (x"f5",x"48",x"73",x"78"),
   241 => (x"5e",x"0e",x"87",x"c8"),
   242 => (x"0e",x"5d",x"5c",x"5b"),
   243 => (x"ff",x"c0",x"1e",x"c0"),
   244 => (x"49",x"c9",x"c1",x"f0"),
   245 => (x"d2",x"87",x"fb",x"f4"),
   246 => (x"e0",x"cd",x"c2",x"1e"),
   247 => (x"87",x"fd",x"fc",x"49"),
   248 => (x"4c",x"c0",x"86",x"c8"),
   249 => (x"b7",x"d2",x"84",x"c1"),
   250 => (x"87",x"f8",x"04",x"ac"),
   251 => (x"97",x"e0",x"cd",x"c2"),
   252 => (x"c0",x"c3",x"49",x"bf"),
   253 => (x"a9",x"c0",x"c1",x"99"),
   254 => (x"87",x"e7",x"c0",x"05"),
   255 => (x"97",x"e7",x"cd",x"c2"),
   256 => (x"31",x"d0",x"49",x"bf"),
   257 => (x"97",x"e8",x"cd",x"c2"),
   258 => (x"32",x"c8",x"4a",x"bf"),
   259 => (x"cd",x"c2",x"b1",x"72"),
   260 => (x"4a",x"bf",x"97",x"e9"),
   261 => (x"cf",x"4c",x"71",x"b1"),
   262 => (x"9c",x"ff",x"ff",x"ff"),
   263 => (x"34",x"ca",x"84",x"c1"),
   264 => (x"c2",x"87",x"e7",x"c1"),
   265 => (x"bf",x"97",x"e9",x"cd"),
   266 => (x"c6",x"31",x"c1",x"49"),
   267 => (x"ea",x"cd",x"c2",x"99"),
   268 => (x"c7",x"4a",x"bf",x"97"),
   269 => (x"b1",x"72",x"2a",x"b7"),
   270 => (x"97",x"e5",x"cd",x"c2"),
   271 => (x"cf",x"4d",x"4a",x"bf"),
   272 => (x"e6",x"cd",x"c2",x"9d"),
   273 => (x"c3",x"4a",x"bf",x"97"),
   274 => (x"c2",x"32",x"ca",x"9a"),
   275 => (x"bf",x"97",x"e7",x"cd"),
   276 => (x"73",x"33",x"c2",x"4b"),
   277 => (x"e8",x"cd",x"c2",x"b2"),
   278 => (x"c3",x"4b",x"bf",x"97"),
   279 => (x"b7",x"c6",x"9b",x"c0"),
   280 => (x"c2",x"b2",x"73",x"2b"),
   281 => (x"71",x"48",x"c1",x"81"),
   282 => (x"c1",x"49",x"70",x"30"),
   283 => (x"70",x"30",x"75",x"48"),
   284 => (x"c1",x"4c",x"72",x"4d"),
   285 => (x"c8",x"94",x"71",x"84"),
   286 => (x"06",x"ad",x"b7",x"c0"),
   287 => (x"34",x"c1",x"87",x"cc"),
   288 => (x"c0",x"c8",x"2d",x"b7"),
   289 => (x"ff",x"01",x"ad",x"b7"),
   290 => (x"48",x"74",x"87",x"f4"),
   291 => (x"0e",x"87",x"fb",x"f1"),
   292 => (x"5d",x"5c",x"5b",x"5e"),
   293 => (x"c2",x"86",x"f8",x"0e"),
   294 => (x"c0",x"48",x"c6",x"d6"),
   295 => (x"fe",x"cd",x"c2",x"78"),
   296 => (x"fb",x"49",x"c0",x"1e"),
   297 => (x"86",x"c4",x"87",x"de"),
   298 => (x"c5",x"05",x"98",x"70"),
   299 => (x"c9",x"48",x"c0",x"87"),
   300 => (x"4d",x"c0",x"87",x"c0"),
   301 => (x"ed",x"c0",x"7e",x"c1"),
   302 => (x"c2",x"49",x"bf",x"e2"),
   303 => (x"71",x"4a",x"f4",x"ce"),
   304 => (x"e4",x"ee",x"4b",x"c8"),
   305 => (x"05",x"98",x"70",x"87"),
   306 => (x"7e",x"c0",x"87",x"c2"),
   307 => (x"bf",x"de",x"ed",x"c0"),
   308 => (x"d0",x"cf",x"c2",x"49"),
   309 => (x"4b",x"c8",x"71",x"4a"),
   310 => (x"70",x"87",x"ce",x"ee"),
   311 => (x"87",x"c2",x"05",x"98"),
   312 => (x"02",x"6e",x"7e",x"c0"),
   313 => (x"c2",x"87",x"fd",x"c0"),
   314 => (x"4d",x"bf",x"c4",x"d5"),
   315 => (x"9f",x"fc",x"d5",x"c2"),
   316 => (x"c5",x"48",x"7e",x"bf"),
   317 => (x"05",x"a8",x"ea",x"d6"),
   318 => (x"d5",x"c2",x"87",x"c7"),
   319 => (x"ce",x"4d",x"bf",x"c4"),
   320 => (x"ca",x"48",x"6e",x"87"),
   321 => (x"02",x"a8",x"d5",x"e9"),
   322 => (x"48",x"c0",x"87",x"c5"),
   323 => (x"c2",x"87",x"e3",x"c7"),
   324 => (x"75",x"1e",x"fe",x"cd"),
   325 => (x"87",x"ec",x"f9",x"49"),
   326 => (x"98",x"70",x"86",x"c4"),
   327 => (x"c0",x"87",x"c5",x"05"),
   328 => (x"87",x"ce",x"c7",x"48"),
   329 => (x"bf",x"de",x"ed",x"c0"),
   330 => (x"d0",x"cf",x"c2",x"49"),
   331 => (x"4b",x"c8",x"71",x"4a"),
   332 => (x"70",x"87",x"f6",x"ec"),
   333 => (x"87",x"c8",x"05",x"98"),
   334 => (x"48",x"c6",x"d6",x"c2"),
   335 => (x"87",x"da",x"78",x"c1"),
   336 => (x"bf",x"e2",x"ed",x"c0"),
   337 => (x"f4",x"ce",x"c2",x"49"),
   338 => (x"4b",x"c8",x"71",x"4a"),
   339 => (x"70",x"87",x"da",x"ec"),
   340 => (x"c5",x"c0",x"02",x"98"),
   341 => (x"c6",x"48",x"c0",x"87"),
   342 => (x"d5",x"c2",x"87",x"d8"),
   343 => (x"49",x"bf",x"97",x"fc"),
   344 => (x"05",x"a9",x"d5",x"c1"),
   345 => (x"c2",x"87",x"cd",x"c0"),
   346 => (x"bf",x"97",x"fd",x"d5"),
   347 => (x"a9",x"ea",x"c2",x"49"),
   348 => (x"87",x"c5",x"c0",x"02"),
   349 => (x"f9",x"c5",x"48",x"c0"),
   350 => (x"fe",x"cd",x"c2",x"87"),
   351 => (x"48",x"7e",x"bf",x"97"),
   352 => (x"02",x"a8",x"e9",x"c3"),
   353 => (x"6e",x"87",x"ce",x"c0"),
   354 => (x"a8",x"eb",x"c3",x"48"),
   355 => (x"87",x"c5",x"c0",x"02"),
   356 => (x"dd",x"c5",x"48",x"c0"),
   357 => (x"c9",x"ce",x"c2",x"87"),
   358 => (x"99",x"49",x"bf",x"97"),
   359 => (x"87",x"cc",x"c0",x"05"),
   360 => (x"97",x"ca",x"ce",x"c2"),
   361 => (x"a9",x"c2",x"49",x"bf"),
   362 => (x"87",x"c5",x"c0",x"02"),
   363 => (x"c1",x"c5",x"48",x"c0"),
   364 => (x"cb",x"ce",x"c2",x"87"),
   365 => (x"c2",x"48",x"bf",x"97"),
   366 => (x"70",x"58",x"c2",x"d6"),
   367 => (x"88",x"c1",x"48",x"4c"),
   368 => (x"58",x"c6",x"d6",x"c2"),
   369 => (x"97",x"cc",x"ce",x"c2"),
   370 => (x"81",x"75",x"49",x"bf"),
   371 => (x"97",x"cd",x"ce",x"c2"),
   372 => (x"32",x"c8",x"4a",x"bf"),
   373 => (x"c2",x"7e",x"a1",x"72"),
   374 => (x"6e",x"48",x"d3",x"da"),
   375 => (x"ce",x"ce",x"c2",x"78"),
   376 => (x"c8",x"48",x"bf",x"97"),
   377 => (x"d6",x"c2",x"58",x"a6"),
   378 => (x"c2",x"02",x"bf",x"c6"),
   379 => (x"ed",x"c0",x"87",x"cf"),
   380 => (x"c2",x"49",x"bf",x"de"),
   381 => (x"71",x"4a",x"d0",x"cf"),
   382 => (x"ec",x"e9",x"4b",x"c8"),
   383 => (x"02",x"98",x"70",x"87"),
   384 => (x"c0",x"87",x"c5",x"c0"),
   385 => (x"87",x"ea",x"c3",x"48"),
   386 => (x"bf",x"fe",x"d5",x"c2"),
   387 => (x"e7",x"da",x"c2",x"4c"),
   388 => (x"e3",x"ce",x"c2",x"5c"),
   389 => (x"c8",x"49",x"bf",x"97"),
   390 => (x"e2",x"ce",x"c2",x"31"),
   391 => (x"a1",x"4a",x"bf",x"97"),
   392 => (x"e4",x"ce",x"c2",x"49"),
   393 => (x"d0",x"4a",x"bf",x"97"),
   394 => (x"49",x"a1",x"72",x"32"),
   395 => (x"97",x"e5",x"ce",x"c2"),
   396 => (x"32",x"d8",x"4a",x"bf"),
   397 => (x"c4",x"49",x"a1",x"72"),
   398 => (x"da",x"c2",x"91",x"66"),
   399 => (x"c2",x"81",x"bf",x"d3"),
   400 => (x"c2",x"59",x"db",x"da"),
   401 => (x"bf",x"97",x"eb",x"ce"),
   402 => (x"c2",x"32",x"c8",x"4a"),
   403 => (x"bf",x"97",x"ea",x"ce"),
   404 => (x"c2",x"4a",x"a2",x"4b"),
   405 => (x"bf",x"97",x"ec",x"ce"),
   406 => (x"73",x"33",x"d0",x"4b"),
   407 => (x"ce",x"c2",x"4a",x"a2"),
   408 => (x"4b",x"bf",x"97",x"ed"),
   409 => (x"33",x"d8",x"9b",x"cf"),
   410 => (x"c2",x"4a",x"a2",x"73"),
   411 => (x"c2",x"5a",x"df",x"da"),
   412 => (x"c2",x"92",x"74",x"8a"),
   413 => (x"72",x"48",x"df",x"da"),
   414 => (x"c1",x"c1",x"78",x"a1"),
   415 => (x"d0",x"ce",x"c2",x"87"),
   416 => (x"c8",x"49",x"bf",x"97"),
   417 => (x"cf",x"ce",x"c2",x"31"),
   418 => (x"a1",x"4a",x"bf",x"97"),
   419 => (x"c7",x"31",x"c5",x"49"),
   420 => (x"29",x"c9",x"81",x"ff"),
   421 => (x"59",x"e7",x"da",x"c2"),
   422 => (x"97",x"d5",x"ce",x"c2"),
   423 => (x"32",x"c8",x"4a",x"bf"),
   424 => (x"97",x"d4",x"ce",x"c2"),
   425 => (x"4a",x"a2",x"4b",x"bf"),
   426 => (x"6e",x"92",x"66",x"c4"),
   427 => (x"e3",x"da",x"c2",x"82"),
   428 => (x"db",x"da",x"c2",x"5a"),
   429 => (x"c2",x"78",x"c0",x"48"),
   430 => (x"72",x"48",x"d7",x"da"),
   431 => (x"da",x"c2",x"78",x"a1"),
   432 => (x"da",x"c2",x"48",x"e7"),
   433 => (x"c2",x"78",x"bf",x"db"),
   434 => (x"c2",x"48",x"eb",x"da"),
   435 => (x"78",x"bf",x"df",x"da"),
   436 => (x"bf",x"c6",x"d6",x"c2"),
   437 => (x"87",x"c9",x"c0",x"02"),
   438 => (x"30",x"c4",x"48",x"74"),
   439 => (x"c9",x"c0",x"7e",x"70"),
   440 => (x"e3",x"da",x"c2",x"87"),
   441 => (x"30",x"c4",x"48",x"bf"),
   442 => (x"d6",x"c2",x"7e",x"70"),
   443 => (x"78",x"6e",x"48",x"ca"),
   444 => (x"8e",x"f8",x"48",x"c1"),
   445 => (x"4c",x"26",x"4d",x"26"),
   446 => (x"4f",x"26",x"4b",x"26"),
   447 => (x"5c",x"5b",x"5e",x"0e"),
   448 => (x"4a",x"71",x"0e",x"5d"),
   449 => (x"bf",x"c6",x"d6",x"c2"),
   450 => (x"72",x"87",x"cb",x"02"),
   451 => (x"72",x"2b",x"c7",x"4b"),
   452 => (x"9d",x"ff",x"c1",x"4d"),
   453 => (x"4b",x"72",x"87",x"c9"),
   454 => (x"4d",x"72",x"2b",x"c8"),
   455 => (x"c2",x"9d",x"ff",x"c3"),
   456 => (x"83",x"bf",x"d3",x"da"),
   457 => (x"bf",x"da",x"ed",x"c0"),
   458 => (x"87",x"d9",x"02",x"ab"),
   459 => (x"5b",x"de",x"ed",x"c0"),
   460 => (x"1e",x"fe",x"cd",x"c2"),
   461 => (x"cb",x"f1",x"49",x"73"),
   462 => (x"70",x"86",x"c4",x"87"),
   463 => (x"87",x"c5",x"05",x"98"),
   464 => (x"e6",x"c0",x"48",x"c0"),
   465 => (x"c6",x"d6",x"c2",x"87"),
   466 => (x"87",x"d2",x"02",x"bf"),
   467 => (x"91",x"c4",x"49",x"75"),
   468 => (x"81",x"fe",x"cd",x"c2"),
   469 => (x"ff",x"cf",x"4c",x"69"),
   470 => (x"9c",x"ff",x"ff",x"ff"),
   471 => (x"49",x"75",x"87",x"cb"),
   472 => (x"cd",x"c2",x"91",x"c2"),
   473 => (x"69",x"9f",x"81",x"fe"),
   474 => (x"fe",x"48",x"74",x"4c"),
   475 => (x"5e",x"0e",x"87",x"c6"),
   476 => (x"0e",x"5d",x"5c",x"5b"),
   477 => (x"4c",x"71",x"86",x"f8"),
   478 => (x"87",x"c5",x"05",x"9c"),
   479 => (x"c0",x"c3",x"48",x"c0"),
   480 => (x"7e",x"a4",x"c8",x"87"),
   481 => (x"d8",x"78",x"c0",x"48"),
   482 => (x"87",x"c7",x"02",x"66"),
   483 => (x"bf",x"97",x"66",x"d8"),
   484 => (x"c0",x"87",x"c5",x"05"),
   485 => (x"87",x"e9",x"c2",x"48"),
   486 => (x"49",x"c1",x"1e",x"c0"),
   487 => (x"87",x"e3",x"c7",x"49"),
   488 => (x"4d",x"70",x"86",x"c4"),
   489 => (x"c2",x"c1",x"02",x"9d"),
   490 => (x"ce",x"d6",x"c2",x"87"),
   491 => (x"49",x"66",x"d8",x"4a"),
   492 => (x"70",x"87",x"db",x"e2"),
   493 => (x"f2",x"c0",x"02",x"98"),
   494 => (x"d8",x"4a",x"75",x"87"),
   495 => (x"4b",x"cb",x"49",x"66"),
   496 => (x"70",x"87",x"c0",x"e3"),
   497 => (x"e2",x"c0",x"02",x"98"),
   498 => (x"75",x"1e",x"c0",x"87"),
   499 => (x"87",x"c7",x"02",x"9d"),
   500 => (x"c0",x"48",x"a6",x"c8"),
   501 => (x"c8",x"87",x"c5",x"78"),
   502 => (x"78",x"c1",x"48",x"a6"),
   503 => (x"c6",x"49",x"66",x"c8"),
   504 => (x"86",x"c4",x"87",x"e1"),
   505 => (x"05",x"9d",x"4d",x"70"),
   506 => (x"75",x"87",x"fe",x"fe"),
   507 => (x"ce",x"c1",x"02",x"9d"),
   508 => (x"49",x"a5",x"dc",x"87"),
   509 => (x"78",x"69",x"48",x"6e"),
   510 => (x"c4",x"49",x"a5",x"da"),
   511 => (x"a4",x"c4",x"48",x"a6"),
   512 => (x"48",x"69",x"9f",x"78"),
   513 => (x"78",x"08",x"66",x"c4"),
   514 => (x"bf",x"c6",x"d6",x"c2"),
   515 => (x"d4",x"87",x"d2",x"02"),
   516 => (x"69",x"9f",x"49",x"a5"),
   517 => (x"ff",x"ff",x"c0",x"49"),
   518 => (x"d0",x"48",x"71",x"99"),
   519 => (x"c2",x"7e",x"70",x"30"),
   520 => (x"6e",x"7e",x"c0",x"87"),
   521 => (x"bf",x"66",x"c4",x"48"),
   522 => (x"08",x"66",x"c4",x"80"),
   523 => (x"cc",x"7c",x"c0",x"78"),
   524 => (x"66",x"c4",x"49",x"a4"),
   525 => (x"a4",x"d0",x"79",x"bf"),
   526 => (x"c1",x"79",x"c0",x"49"),
   527 => (x"c0",x"87",x"c2",x"48"),
   528 => (x"fa",x"8e",x"f8",x"48"),
   529 => (x"5e",x"0e",x"87",x"ee"),
   530 => (x"71",x"0e",x"5c",x"5b"),
   531 => (x"c1",x"02",x"9c",x"4c"),
   532 => (x"a4",x"c8",x"87",x"cb"),
   533 => (x"c1",x"02",x"69",x"49"),
   534 => (x"49",x"6c",x"87",x"c3"),
   535 => (x"71",x"48",x"66",x"cc"),
   536 => (x"58",x"a6",x"d0",x"80"),
   537 => (x"d6",x"c2",x"b9",x"70"),
   538 => (x"ff",x"4a",x"bf",x"c2"),
   539 => (x"71",x"99",x"72",x"ba"),
   540 => (x"e5",x"c0",x"02",x"99"),
   541 => (x"4b",x"a4",x"c4",x"87"),
   542 => (x"ff",x"f9",x"49",x"6b"),
   543 => (x"c2",x"7b",x"70",x"87"),
   544 => (x"49",x"bf",x"fe",x"d5"),
   545 => (x"7c",x"71",x"81",x"6c"),
   546 => (x"c2",x"b9",x"66",x"cc"),
   547 => (x"4a",x"bf",x"c2",x"d6"),
   548 => (x"99",x"72",x"ba",x"ff"),
   549 => (x"ff",x"05",x"99",x"71"),
   550 => (x"66",x"cc",x"87",x"db"),
   551 => (x"87",x"d6",x"f9",x"7c"),
   552 => (x"71",x"1e",x"73",x"1e"),
   553 => (x"c7",x"02",x"9b",x"4b"),
   554 => (x"49",x"a3",x"c8",x"87"),
   555 => (x"87",x"c5",x"05",x"69"),
   556 => (x"f6",x"c0",x"48",x"c0"),
   557 => (x"d7",x"da",x"c2",x"87"),
   558 => (x"a3",x"c4",x"49",x"bf"),
   559 => (x"c2",x"4a",x"6a",x"4a"),
   560 => (x"fe",x"d5",x"c2",x"8a"),
   561 => (x"a1",x"72",x"92",x"bf"),
   562 => (x"c2",x"d6",x"c2",x"49"),
   563 => (x"9a",x"6b",x"4a",x"bf"),
   564 => (x"c0",x"49",x"a1",x"72"),
   565 => (x"c8",x"59",x"de",x"ed"),
   566 => (x"ea",x"71",x"1e",x"66"),
   567 => (x"86",x"c4",x"87",x"e6"),
   568 => (x"c4",x"05",x"98",x"70"),
   569 => (x"c2",x"48",x"c0",x"87"),
   570 => (x"f8",x"48",x"c1",x"87"),
   571 => (x"73",x"1e",x"87",x"ca"),
   572 => (x"9b",x"4b",x"71",x"1e"),
   573 => (x"87",x"e4",x"c0",x"02"),
   574 => (x"5b",x"eb",x"da",x"c2"),
   575 => (x"8a",x"c2",x"4a",x"73"),
   576 => (x"bf",x"fe",x"d5",x"c2"),
   577 => (x"da",x"c2",x"92",x"49"),
   578 => (x"72",x"48",x"bf",x"d7"),
   579 => (x"ef",x"da",x"c2",x"80"),
   580 => (x"c4",x"48",x"71",x"58"),
   581 => (x"ce",x"d6",x"c2",x"30"),
   582 => (x"87",x"ed",x"c0",x"58"),
   583 => (x"48",x"e7",x"da",x"c2"),
   584 => (x"bf",x"db",x"da",x"c2"),
   585 => (x"eb",x"da",x"c2",x"78"),
   586 => (x"df",x"da",x"c2",x"48"),
   587 => (x"d6",x"c2",x"78",x"bf"),
   588 => (x"c9",x"02",x"bf",x"c6"),
   589 => (x"fe",x"d5",x"c2",x"87"),
   590 => (x"31",x"c4",x"49",x"bf"),
   591 => (x"da",x"c2",x"87",x"c7"),
   592 => (x"c4",x"49",x"bf",x"e3"),
   593 => (x"ce",x"d6",x"c2",x"31"),
   594 => (x"87",x"ec",x"f6",x"59"),
   595 => (x"5c",x"5b",x"5e",x"0e"),
   596 => (x"c0",x"4a",x"71",x"0e"),
   597 => (x"02",x"9a",x"72",x"4b"),
   598 => (x"da",x"87",x"e0",x"c0"),
   599 => (x"69",x"9f",x"49",x"a2"),
   600 => (x"c6",x"d6",x"c2",x"4b"),
   601 => (x"87",x"cf",x"02",x"bf"),
   602 => (x"9f",x"49",x"a2",x"d4"),
   603 => (x"c0",x"4c",x"49",x"69"),
   604 => (x"d0",x"9c",x"ff",x"ff"),
   605 => (x"c0",x"87",x"c2",x"34"),
   606 => (x"73",x"b3",x"74",x"4c"),
   607 => (x"87",x"ee",x"fd",x"49"),
   608 => (x"0e",x"87",x"f3",x"f5"),
   609 => (x"5d",x"5c",x"5b",x"5e"),
   610 => (x"71",x"86",x"f4",x"0e"),
   611 => (x"72",x"7e",x"c0",x"4a"),
   612 => (x"87",x"d8",x"02",x"9a"),
   613 => (x"48",x"fa",x"cd",x"c2"),
   614 => (x"cd",x"c2",x"78",x"c0"),
   615 => (x"da",x"c2",x"48",x"f2"),
   616 => (x"c2",x"78",x"bf",x"eb"),
   617 => (x"c2",x"48",x"f6",x"cd"),
   618 => (x"78",x"bf",x"e7",x"da"),
   619 => (x"48",x"db",x"d6",x"c2"),
   620 => (x"d6",x"c2",x"50",x"c0"),
   621 => (x"c2",x"49",x"bf",x"ca"),
   622 => (x"4a",x"bf",x"fa",x"cd"),
   623 => (x"c4",x"03",x"aa",x"71"),
   624 => (x"49",x"72",x"87",x"c9"),
   625 => (x"c0",x"05",x"99",x"cf"),
   626 => (x"ed",x"c0",x"87",x"e9"),
   627 => (x"cd",x"c2",x"48",x"da"),
   628 => (x"c2",x"78",x"bf",x"f2"),
   629 => (x"c2",x"1e",x"fe",x"cd"),
   630 => (x"49",x"bf",x"f2",x"cd"),
   631 => (x"48",x"f2",x"cd",x"c2"),
   632 => (x"71",x"78",x"a1",x"c1"),
   633 => (x"c4",x"87",x"dd",x"e6"),
   634 => (x"d6",x"ed",x"c0",x"86"),
   635 => (x"fe",x"cd",x"c2",x"48"),
   636 => (x"c0",x"87",x"cc",x"78"),
   637 => (x"48",x"bf",x"d6",x"ed"),
   638 => (x"c0",x"80",x"e0",x"c0"),
   639 => (x"c2",x"58",x"da",x"ed"),
   640 => (x"48",x"bf",x"fa",x"cd"),
   641 => (x"cd",x"c2",x"80",x"c1"),
   642 => (x"56",x"27",x"58",x"fe"),
   643 => (x"bf",x"00",x"00",x"0b"),
   644 => (x"9d",x"4d",x"bf",x"97"),
   645 => (x"87",x"e3",x"c2",x"02"),
   646 => (x"02",x"ad",x"e5",x"c3"),
   647 => (x"c0",x"87",x"dc",x"c2"),
   648 => (x"4b",x"bf",x"d6",x"ed"),
   649 => (x"11",x"49",x"a3",x"cb"),
   650 => (x"05",x"ac",x"cf",x"4c"),
   651 => (x"75",x"87",x"d2",x"c1"),
   652 => (x"c1",x"99",x"df",x"49"),
   653 => (x"c2",x"91",x"cd",x"89"),
   654 => (x"c1",x"81",x"ce",x"d6"),
   655 => (x"51",x"12",x"4a",x"a3"),
   656 => (x"12",x"4a",x"a3",x"c3"),
   657 => (x"4a",x"a3",x"c5",x"51"),
   658 => (x"a3",x"c7",x"51",x"12"),
   659 => (x"c9",x"51",x"12",x"4a"),
   660 => (x"51",x"12",x"4a",x"a3"),
   661 => (x"12",x"4a",x"a3",x"ce"),
   662 => (x"4a",x"a3",x"d0",x"51"),
   663 => (x"a3",x"d2",x"51",x"12"),
   664 => (x"d4",x"51",x"12",x"4a"),
   665 => (x"51",x"12",x"4a",x"a3"),
   666 => (x"12",x"4a",x"a3",x"d6"),
   667 => (x"4a",x"a3",x"d8",x"51"),
   668 => (x"a3",x"dc",x"51",x"12"),
   669 => (x"de",x"51",x"12",x"4a"),
   670 => (x"51",x"12",x"4a",x"a3"),
   671 => (x"fa",x"c0",x"7e",x"c1"),
   672 => (x"c8",x"49",x"74",x"87"),
   673 => (x"eb",x"c0",x"05",x"99"),
   674 => (x"d0",x"49",x"74",x"87"),
   675 => (x"87",x"d1",x"05",x"99"),
   676 => (x"c0",x"02",x"66",x"dc"),
   677 => (x"49",x"73",x"87",x"cb"),
   678 => (x"70",x"0f",x"66",x"dc"),
   679 => (x"d3",x"c0",x"02",x"98"),
   680 => (x"c0",x"05",x"6e",x"87"),
   681 => (x"d6",x"c2",x"87",x"c6"),
   682 => (x"50",x"c0",x"48",x"ce"),
   683 => (x"bf",x"d6",x"ed",x"c0"),
   684 => (x"87",x"dd",x"c2",x"48"),
   685 => (x"48",x"db",x"d6",x"c2"),
   686 => (x"c2",x"7e",x"50",x"c0"),
   687 => (x"49",x"bf",x"ca",x"d6"),
   688 => (x"bf",x"fa",x"cd",x"c2"),
   689 => (x"04",x"aa",x"71",x"4a"),
   690 => (x"c2",x"87",x"f7",x"fb"),
   691 => (x"05",x"bf",x"eb",x"da"),
   692 => (x"c2",x"87",x"c8",x"c0"),
   693 => (x"02",x"bf",x"c6",x"d6"),
   694 => (x"c2",x"87",x"f4",x"c1"),
   695 => (x"49",x"bf",x"f6",x"cd"),
   696 => (x"c2",x"87",x"d9",x"f0"),
   697 => (x"c4",x"58",x"fa",x"cd"),
   698 => (x"cd",x"c2",x"48",x"a6"),
   699 => (x"c2",x"78",x"bf",x"f6"),
   700 => (x"02",x"bf",x"c6",x"d6"),
   701 => (x"c4",x"87",x"d8",x"c0"),
   702 => (x"ff",x"cf",x"49",x"66"),
   703 => (x"99",x"f8",x"ff",x"ff"),
   704 => (x"c5",x"c0",x"02",x"a9"),
   705 => (x"c0",x"4c",x"c0",x"87"),
   706 => (x"4c",x"c1",x"87",x"e1"),
   707 => (x"c4",x"87",x"dc",x"c0"),
   708 => (x"ff",x"cf",x"49",x"66"),
   709 => (x"02",x"a9",x"99",x"f8"),
   710 => (x"c8",x"87",x"c8",x"c0"),
   711 => (x"78",x"c0",x"48",x"a6"),
   712 => (x"c8",x"87",x"c5",x"c0"),
   713 => (x"78",x"c1",x"48",x"a6"),
   714 => (x"74",x"4c",x"66",x"c8"),
   715 => (x"de",x"c0",x"05",x"9c"),
   716 => (x"49",x"66",x"c4",x"87"),
   717 => (x"d5",x"c2",x"89",x"c2"),
   718 => (x"c2",x"91",x"bf",x"fe"),
   719 => (x"48",x"bf",x"d7",x"da"),
   720 => (x"cd",x"c2",x"80",x"71"),
   721 => (x"cd",x"c2",x"58",x"f6"),
   722 => (x"78",x"c0",x"48",x"fa"),
   723 => (x"c0",x"87",x"e3",x"f9"),
   724 => (x"ee",x"8e",x"f4",x"48"),
   725 => (x"00",x"00",x"87",x"de"),
   726 => (x"ff",x"ff",x"00",x"00"),
   727 => (x"0b",x"66",x"ff",x"ff"),
   728 => (x"0b",x"6f",x"00",x"00"),
   729 => (x"41",x"46",x"00",x"00"),
   730 => (x"20",x"32",x"33",x"54"),
   731 => (x"46",x"00",x"20",x"20"),
   732 => (x"36",x"31",x"54",x"41"),
   733 => (x"00",x"20",x"20",x"20"),
   734 => (x"48",x"d4",x"ff",x"1e"),
   735 => (x"68",x"78",x"ff",x"c3"),
   736 => (x"1e",x"4f",x"26",x"48"),
   737 => (x"c3",x"48",x"d4",x"ff"),
   738 => (x"d0",x"ff",x"78",x"ff"),
   739 => (x"78",x"e1",x"c0",x"48"),
   740 => (x"d4",x"48",x"d4",x"ff"),
   741 => (x"ef",x"da",x"c2",x"78"),
   742 => (x"bf",x"d4",x"ff",x"48"),
   743 => (x"1e",x"4f",x"26",x"50"),
   744 => (x"c0",x"48",x"d0",x"ff"),
   745 => (x"4f",x"26",x"78",x"e0"),
   746 => (x"87",x"cc",x"ff",x"1e"),
   747 => (x"02",x"99",x"49",x"70"),
   748 => (x"fb",x"c0",x"87",x"c6"),
   749 => (x"87",x"f1",x"05",x"a9"),
   750 => (x"4f",x"26",x"48",x"71"),
   751 => (x"5c",x"5b",x"5e",x"0e"),
   752 => (x"c0",x"4b",x"71",x"0e"),
   753 => (x"87",x"f0",x"fe",x"4c"),
   754 => (x"02",x"99",x"49",x"70"),
   755 => (x"c0",x"87",x"f9",x"c0"),
   756 => (x"c0",x"02",x"a9",x"ec"),
   757 => (x"fb",x"c0",x"87",x"f2"),
   758 => (x"eb",x"c0",x"02",x"a9"),
   759 => (x"b7",x"66",x"cc",x"87"),
   760 => (x"87",x"c7",x"03",x"ac"),
   761 => (x"c2",x"02",x"66",x"d0"),
   762 => (x"71",x"53",x"71",x"87"),
   763 => (x"87",x"c2",x"02",x"99"),
   764 => (x"c3",x"fe",x"84",x"c1"),
   765 => (x"99",x"49",x"70",x"87"),
   766 => (x"c0",x"87",x"cd",x"02"),
   767 => (x"c7",x"02",x"a9",x"ec"),
   768 => (x"a9",x"fb",x"c0",x"87"),
   769 => (x"87",x"d5",x"ff",x"05"),
   770 => (x"c3",x"02",x"66",x"d0"),
   771 => (x"7b",x"97",x"c0",x"87"),
   772 => (x"05",x"a9",x"ec",x"c0"),
   773 => (x"4a",x"74",x"87",x"c4"),
   774 => (x"4a",x"74",x"87",x"c5"),
   775 => (x"72",x"8a",x"0a",x"c0"),
   776 => (x"26",x"87",x"c2",x"48"),
   777 => (x"26",x"4c",x"26",x"4d"),
   778 => (x"1e",x"4f",x"26",x"4b"),
   779 => (x"70",x"87",x"c9",x"fd"),
   780 => (x"f0",x"c0",x"4a",x"49"),
   781 => (x"87",x"c9",x"04",x"aa"),
   782 => (x"01",x"aa",x"f9",x"c0"),
   783 => (x"f0",x"c0",x"87",x"c3"),
   784 => (x"aa",x"c1",x"c1",x"8a"),
   785 => (x"c1",x"87",x"c9",x"04"),
   786 => (x"c3",x"01",x"aa",x"da"),
   787 => (x"8a",x"f7",x"c0",x"87"),
   788 => (x"4f",x"26",x"48",x"72"),
   789 => (x"5c",x"5b",x"5e",x"0e"),
   790 => (x"86",x"f8",x"0e",x"5d"),
   791 => (x"4d",x"c0",x"4c",x"71"),
   792 => (x"c0",x"87",x"e0",x"fc"),
   793 => (x"f3",x"f3",x"c0",x"4b"),
   794 => (x"c0",x"49",x"bf",x"97"),
   795 => (x"87",x"cf",x"04",x"a9"),
   796 => (x"c1",x"87",x"f5",x"fc"),
   797 => (x"f3",x"f3",x"c0",x"83"),
   798 => (x"ab",x"49",x"bf",x"97"),
   799 => (x"c0",x"87",x"f1",x"06"),
   800 => (x"bf",x"97",x"f3",x"f3"),
   801 => (x"fb",x"87",x"cf",x"02"),
   802 => (x"49",x"70",x"87",x"ee"),
   803 => (x"87",x"c6",x"02",x"99"),
   804 => (x"05",x"a9",x"ec",x"c0"),
   805 => (x"4b",x"c0",x"87",x"f1"),
   806 => (x"70",x"87",x"dd",x"fb"),
   807 => (x"87",x"d8",x"fb",x"7e"),
   808 => (x"fb",x"58",x"a6",x"c8"),
   809 => (x"4a",x"70",x"87",x"d2"),
   810 => (x"a4",x"c8",x"83",x"c1"),
   811 => (x"49",x"69",x"97",x"49"),
   812 => (x"da",x"05",x"a9",x"6e"),
   813 => (x"49",x"a4",x"c9",x"87"),
   814 => (x"c4",x"49",x"69",x"97"),
   815 => (x"ce",x"05",x"a9",x"66"),
   816 => (x"49",x"a4",x"ca",x"87"),
   817 => (x"aa",x"49",x"69",x"97"),
   818 => (x"c1",x"87",x"c4",x"05"),
   819 => (x"6e",x"87",x"d4",x"4d"),
   820 => (x"a8",x"ec",x"c0",x"48"),
   821 => (x"6e",x"87",x"c8",x"02"),
   822 => (x"a8",x"fb",x"c0",x"48"),
   823 => (x"c0",x"87",x"c4",x"05"),
   824 => (x"75",x"4d",x"c1",x"4b"),
   825 => (x"ef",x"fe",x"02",x"9d"),
   826 => (x"87",x"f3",x"fa",x"87"),
   827 => (x"8e",x"f8",x"48",x"73"),
   828 => (x"00",x"87",x"f0",x"fc"),
   829 => (x"5c",x"5b",x"5e",x"0e"),
   830 => (x"86",x"f8",x"0e",x"5d"),
   831 => (x"d4",x"ff",x"7e",x"71"),
   832 => (x"c2",x"1e",x"6e",x"4b"),
   833 => (x"e9",x"49",x"f4",x"da"),
   834 => (x"86",x"c4",x"87",x"e4"),
   835 => (x"c4",x"02",x"98",x"70"),
   836 => (x"dd",x"c1",x"87",x"ea"),
   837 => (x"6e",x"4d",x"bf",x"ec"),
   838 => (x"87",x"f8",x"fc",x"49"),
   839 => (x"70",x"58",x"a6",x"c8"),
   840 => (x"87",x"c5",x"05",x"98"),
   841 => (x"c1",x"48",x"a6",x"c4"),
   842 => (x"48",x"d0",x"ff",x"78"),
   843 => (x"d5",x"c1",x"78",x"c5"),
   844 => (x"49",x"66",x"c4",x"7b"),
   845 => (x"31",x"c6",x"89",x"c1"),
   846 => (x"97",x"ea",x"dd",x"c1"),
   847 => (x"71",x"48",x"4a",x"bf"),
   848 => (x"ff",x"7b",x"70",x"b0"),
   849 => (x"78",x"c4",x"48",x"d0"),
   850 => (x"97",x"ef",x"da",x"c2"),
   851 => (x"99",x"d0",x"49",x"bf"),
   852 => (x"c5",x"87",x"d7",x"02"),
   853 => (x"7b",x"d6",x"c1",x"78"),
   854 => (x"ff",x"c3",x"4a",x"c0"),
   855 => (x"c0",x"82",x"c1",x"7b"),
   856 => (x"f5",x"04",x"aa",x"e0"),
   857 => (x"48",x"d0",x"ff",x"87"),
   858 => (x"ff",x"c3",x"78",x"c4"),
   859 => (x"48",x"d0",x"ff",x"7b"),
   860 => (x"d3",x"c1",x"78",x"c5"),
   861 => (x"c4",x"7b",x"c1",x"7b"),
   862 => (x"ad",x"b7",x"c0",x"78"),
   863 => (x"87",x"eb",x"c2",x"06"),
   864 => (x"bf",x"fc",x"da",x"c2"),
   865 => (x"02",x"9c",x"8d",x"4c"),
   866 => (x"c2",x"87",x"c2",x"c2"),
   867 => (x"c4",x"7e",x"fe",x"cd"),
   868 => (x"c0",x"c8",x"48",x"a6"),
   869 => (x"b7",x"c0",x"8c",x"78"),
   870 => (x"87",x"c6",x"03",x"ac"),
   871 => (x"78",x"a4",x"c0",x"c8"),
   872 => (x"da",x"c2",x"4c",x"c0"),
   873 => (x"49",x"bf",x"97",x"ef"),
   874 => (x"d0",x"02",x"99",x"d0"),
   875 => (x"c2",x"1e",x"c0",x"87"),
   876 => (x"eb",x"49",x"f4",x"da"),
   877 => (x"86",x"c4",x"87",x"ea"),
   878 => (x"f5",x"c0",x"4a",x"70"),
   879 => (x"fe",x"cd",x"c2",x"87"),
   880 => (x"f4",x"da",x"c2",x"1e"),
   881 => (x"87",x"d8",x"eb",x"49"),
   882 => (x"4a",x"70",x"86",x"c4"),
   883 => (x"c8",x"48",x"d0",x"ff"),
   884 => (x"d4",x"c1",x"78",x"c5"),
   885 => (x"bf",x"97",x"6e",x"7b"),
   886 => (x"c1",x"48",x"6e",x"7b"),
   887 => (x"c4",x"7e",x"70",x"80"),
   888 => (x"88",x"c1",x"48",x"66"),
   889 => (x"70",x"58",x"a6",x"c8"),
   890 => (x"e8",x"ff",x"05",x"98"),
   891 => (x"48",x"d0",x"ff",x"87"),
   892 => (x"9a",x"72",x"78",x"c4"),
   893 => (x"c0",x"87",x"c5",x"05"),
   894 => (x"87",x"c2",x"c1",x"48"),
   895 => (x"da",x"c2",x"1e",x"c1"),
   896 => (x"c1",x"e9",x"49",x"f4"),
   897 => (x"74",x"86",x"c4",x"87"),
   898 => (x"fe",x"fd",x"05",x"9c"),
   899 => (x"ad",x"b7",x"c0",x"87"),
   900 => (x"c2",x"87",x"d1",x"06"),
   901 => (x"c0",x"48",x"f4",x"da"),
   902 => (x"c0",x"80",x"d0",x"78"),
   903 => (x"c2",x"80",x"f4",x"78"),
   904 => (x"78",x"bf",x"c0",x"db"),
   905 => (x"01",x"ad",x"b7",x"c0"),
   906 => (x"ff",x"87",x"d5",x"fd"),
   907 => (x"78",x"c5",x"48",x"d0"),
   908 => (x"c0",x"7b",x"d3",x"c1"),
   909 => (x"c1",x"78",x"c4",x"7b"),
   910 => (x"87",x"c2",x"c0",x"48"),
   911 => (x"8e",x"f8",x"48",x"c0"),
   912 => (x"4c",x"26",x"4d",x"26"),
   913 => (x"4f",x"26",x"4b",x"26"),
   914 => (x"5c",x"5b",x"5e",x"0e"),
   915 => (x"71",x"1e",x"0e",x"5d"),
   916 => (x"4d",x"4c",x"c0",x"4b"),
   917 => (x"e8",x"c0",x"04",x"ab"),
   918 => (x"d4",x"f1",x"c0",x"87"),
   919 => (x"02",x"9d",x"75",x"1e"),
   920 => (x"4a",x"c0",x"87",x"c4"),
   921 => (x"4a",x"c1",x"87",x"c2"),
   922 => (x"d6",x"ec",x"49",x"72"),
   923 => (x"70",x"86",x"c4",x"87"),
   924 => (x"6e",x"84",x"c1",x"7e"),
   925 => (x"73",x"87",x"c2",x"05"),
   926 => (x"73",x"85",x"c1",x"4c"),
   927 => (x"d8",x"ff",x"06",x"ac"),
   928 => (x"26",x"48",x"6e",x"87"),
   929 => (x"1e",x"87",x"f9",x"fe"),
   930 => (x"66",x"c4",x"4a",x"71"),
   931 => (x"72",x"87",x"c5",x"05"),
   932 => (x"87",x"e0",x"f9",x"49"),
   933 => (x"5e",x"0e",x"4f",x"26"),
   934 => (x"0e",x"5d",x"5c",x"5b"),
   935 => (x"49",x"4c",x"71",x"1e"),
   936 => (x"db",x"c2",x"91",x"de"),
   937 => (x"85",x"71",x"4d",x"dc"),
   938 => (x"c1",x"02",x"6d",x"97"),
   939 => (x"db",x"c2",x"87",x"dc"),
   940 => (x"74",x"49",x"bf",x"c8"),
   941 => (x"cf",x"fe",x"71",x"81"),
   942 => (x"48",x"7e",x"70",x"87"),
   943 => (x"f2",x"c0",x"02",x"98"),
   944 => (x"d0",x"db",x"c2",x"87"),
   945 => (x"cb",x"4a",x"70",x"4b"),
   946 => (x"da",x"c7",x"ff",x"49"),
   947 => (x"cb",x"4b",x"74",x"87"),
   948 => (x"fe",x"dd",x"c1",x"93"),
   949 => (x"c0",x"83",x"c4",x"83"),
   950 => (x"74",x"7b",x"ce",x"fc"),
   951 => (x"ea",x"c0",x"c1",x"49"),
   952 => (x"c1",x"7b",x"75",x"87"),
   953 => (x"bf",x"97",x"eb",x"dd"),
   954 => (x"db",x"c2",x"1e",x"49"),
   955 => (x"d6",x"fe",x"49",x"d0"),
   956 => (x"74",x"86",x"c4",x"87"),
   957 => (x"d2",x"c0",x"c1",x"49"),
   958 => (x"c1",x"49",x"c0",x"87"),
   959 => (x"c2",x"87",x"f1",x"c1"),
   960 => (x"c0",x"48",x"f0",x"da"),
   961 => (x"de",x"49",x"c1",x"78"),
   962 => (x"fc",x"26",x"87",x"cb"),
   963 => (x"6f",x"4c",x"87",x"f2"),
   964 => (x"6e",x"69",x"64",x"61"),
   965 => (x"2e",x"2e",x"2e",x"67"),
   966 => (x"1e",x"73",x"1e",x"00"),
   967 => (x"c2",x"49",x"4a",x"71"),
   968 => (x"81",x"bf",x"c8",x"db"),
   969 => (x"87",x"e0",x"fc",x"71"),
   970 => (x"02",x"9b",x"4b",x"70"),
   971 => (x"e8",x"49",x"87",x"c4"),
   972 => (x"db",x"c2",x"87",x"da"),
   973 => (x"78",x"c0",x"48",x"c8"),
   974 => (x"d8",x"dd",x"49",x"c1"),
   975 => (x"87",x"c4",x"fc",x"87"),
   976 => (x"c1",x"49",x"c0",x"1e"),
   977 => (x"26",x"87",x"e9",x"c0"),
   978 => (x"4a",x"71",x"1e",x"4f"),
   979 => (x"c1",x"91",x"cb",x"49"),
   980 => (x"c8",x"81",x"fe",x"dd"),
   981 => (x"c2",x"48",x"11",x"81"),
   982 => (x"c2",x"58",x"f4",x"da"),
   983 => (x"c0",x"48",x"c8",x"db"),
   984 => (x"dc",x"49",x"c1",x"78"),
   985 => (x"4f",x"26",x"87",x"ef"),
   986 => (x"02",x"99",x"71",x"1e"),
   987 => (x"df",x"c1",x"87",x"d2"),
   988 => (x"50",x"c0",x"48",x"d3"),
   989 => (x"fd",x"c0",x"80",x"f7"),
   990 => (x"dd",x"c1",x"40",x"c9"),
   991 => (x"87",x"ce",x"78",x"f7"),
   992 => (x"48",x"cf",x"df",x"c1"),
   993 => (x"78",x"f0",x"dd",x"c1"),
   994 => (x"fd",x"c0",x"80",x"fc"),
   995 => (x"4f",x"26",x"78",x"c0"),
   996 => (x"5c",x"5b",x"5e",x"0e"),
   997 => (x"86",x"f4",x"0e",x"5d"),
   998 => (x"4d",x"fe",x"cd",x"c2"),
   999 => (x"a6",x"c4",x"4c",x"c0"),
  1000 => (x"c2",x"78",x"c0",x"48"),
  1001 => (x"48",x"bf",x"c8",x"db"),
  1002 => (x"c1",x"06",x"a8",x"c0"),
  1003 => (x"cd",x"c2",x"87",x"c0"),
  1004 => (x"02",x"98",x"48",x"fe"),
  1005 => (x"c0",x"87",x"f7",x"c0"),
  1006 => (x"c8",x"1e",x"d4",x"f1"),
  1007 => (x"87",x"c7",x"02",x"66"),
  1008 => (x"c0",x"48",x"a6",x"c4"),
  1009 => (x"c4",x"87",x"c5",x"78"),
  1010 => (x"78",x"c1",x"48",x"a6"),
  1011 => (x"e6",x"49",x"66",x"c4"),
  1012 => (x"86",x"c4",x"87",x"f1"),
  1013 => (x"84",x"c1",x"4d",x"70"),
  1014 => (x"c1",x"48",x"66",x"c4"),
  1015 => (x"58",x"a6",x"c8",x"80"),
  1016 => (x"bf",x"c8",x"db",x"c2"),
  1017 => (x"87",x"c6",x"03",x"ac"),
  1018 => (x"ff",x"05",x"9d",x"75"),
  1019 => (x"4c",x"c0",x"87",x"c9"),
  1020 => (x"c3",x"02",x"9d",x"75"),
  1021 => (x"f1",x"c0",x"87",x"dc"),
  1022 => (x"66",x"c8",x"1e",x"d4"),
  1023 => (x"cc",x"87",x"c7",x"02"),
  1024 => (x"78",x"c0",x"48",x"a6"),
  1025 => (x"a6",x"cc",x"87",x"c5"),
  1026 => (x"cc",x"78",x"c1",x"48"),
  1027 => (x"f2",x"e5",x"49",x"66"),
  1028 => (x"70",x"86",x"c4",x"87"),
  1029 => (x"02",x"98",x"48",x"7e"),
  1030 => (x"49",x"87",x"e4",x"c2"),
  1031 => (x"69",x"97",x"81",x"cb"),
  1032 => (x"02",x"99",x"d0",x"49"),
  1033 => (x"74",x"87",x"d4",x"c1"),
  1034 => (x"c1",x"91",x"cb",x"49"),
  1035 => (x"c0",x"81",x"fe",x"dd"),
  1036 => (x"c8",x"79",x"d9",x"fc"),
  1037 => (x"51",x"ff",x"c3",x"81"),
  1038 => (x"91",x"de",x"49",x"74"),
  1039 => (x"4d",x"dc",x"db",x"c2"),
  1040 => (x"c1",x"c2",x"85",x"71"),
  1041 => (x"a5",x"c1",x"7d",x"97"),
  1042 => (x"51",x"e0",x"c0",x"49"),
  1043 => (x"97",x"ce",x"d6",x"c2"),
  1044 => (x"87",x"d2",x"02",x"bf"),
  1045 => (x"a5",x"c2",x"84",x"c1"),
  1046 => (x"ce",x"d6",x"c2",x"4b"),
  1047 => (x"ff",x"49",x"db",x"4a"),
  1048 => (x"c1",x"87",x"c4",x"c1"),
  1049 => (x"a5",x"cd",x"87",x"d9"),
  1050 => (x"c1",x"51",x"c0",x"49"),
  1051 => (x"4b",x"a5",x"c2",x"84"),
  1052 => (x"49",x"cb",x"4a",x"6e"),
  1053 => (x"87",x"ef",x"c0",x"ff"),
  1054 => (x"74",x"87",x"c4",x"c1"),
  1055 => (x"c1",x"91",x"cb",x"49"),
  1056 => (x"c0",x"81",x"fe",x"dd"),
  1057 => (x"c2",x"79",x"d6",x"fa"),
  1058 => (x"bf",x"97",x"ce",x"d6"),
  1059 => (x"74",x"87",x"d8",x"02"),
  1060 => (x"c1",x"91",x"de",x"49"),
  1061 => (x"dc",x"db",x"c2",x"84"),
  1062 => (x"c2",x"83",x"71",x"4b"),
  1063 => (x"dd",x"4a",x"ce",x"d6"),
  1064 => (x"c2",x"c0",x"ff",x"49"),
  1065 => (x"74",x"87",x"d8",x"87"),
  1066 => (x"c2",x"93",x"de",x"4b"),
  1067 => (x"cb",x"83",x"dc",x"db"),
  1068 => (x"51",x"c0",x"49",x"a3"),
  1069 => (x"6e",x"73",x"84",x"c1"),
  1070 => (x"fe",x"49",x"cb",x"4a"),
  1071 => (x"c4",x"87",x"e8",x"ff"),
  1072 => (x"80",x"c1",x"48",x"66"),
  1073 => (x"c7",x"58",x"a6",x"c8"),
  1074 => (x"c5",x"c0",x"03",x"ac"),
  1075 => (x"fc",x"05",x"6e",x"87"),
  1076 => (x"48",x"74",x"87",x"e4"),
  1077 => (x"e7",x"f5",x"8e",x"f4"),
  1078 => (x"1e",x"73",x"1e",x"87"),
  1079 => (x"cb",x"49",x"4b",x"71"),
  1080 => (x"fe",x"dd",x"c1",x"91"),
  1081 => (x"4a",x"a1",x"c8",x"81"),
  1082 => (x"48",x"ea",x"dd",x"c1"),
  1083 => (x"a1",x"c9",x"50",x"12"),
  1084 => (x"f3",x"f3",x"c0",x"4a"),
  1085 => (x"ca",x"50",x"12",x"48"),
  1086 => (x"eb",x"dd",x"c1",x"81"),
  1087 => (x"c1",x"50",x"11",x"48"),
  1088 => (x"bf",x"97",x"eb",x"dd"),
  1089 => (x"49",x"c0",x"1e",x"49"),
  1090 => (x"c2",x"87",x"fc",x"f5"),
  1091 => (x"de",x"48",x"f0",x"da"),
  1092 => (x"d5",x"49",x"c1",x"78"),
  1093 => (x"f4",x"26",x"87",x"ff"),
  1094 => (x"5e",x"0e",x"87",x"ea"),
  1095 => (x"0e",x"5d",x"5c",x"5b"),
  1096 => (x"4d",x"71",x"86",x"f4"),
  1097 => (x"c1",x"91",x"cb",x"49"),
  1098 => (x"c8",x"81",x"fe",x"dd"),
  1099 => (x"a1",x"ca",x"4a",x"a1"),
  1100 => (x"48",x"a6",x"c4",x"7e"),
  1101 => (x"bf",x"f8",x"de",x"c2"),
  1102 => (x"bf",x"97",x"6e",x"78"),
  1103 => (x"48",x"66",x"c4",x"4b"),
  1104 => (x"4b",x"70",x"28",x"73"),
  1105 => (x"cc",x"48",x"12",x"4c"),
  1106 => (x"9c",x"70",x"58",x"a6"),
  1107 => (x"81",x"c9",x"84",x"c1"),
  1108 => (x"b7",x"49",x"69",x"97"),
  1109 => (x"87",x"c2",x"04",x"ac"),
  1110 => (x"97",x"6e",x"4c",x"c0"),
  1111 => (x"66",x"c8",x"4a",x"bf"),
  1112 => (x"ff",x"31",x"72",x"49"),
  1113 => (x"99",x"66",x"c4",x"b9"),
  1114 => (x"30",x"72",x"48",x"74"),
  1115 => (x"71",x"48",x"4a",x"70"),
  1116 => (x"fc",x"de",x"c2",x"b0"),
  1117 => (x"d2",x"e4",x"c0",x"58"),
  1118 => (x"d4",x"49",x"c0",x"87"),
  1119 => (x"49",x"75",x"87",x"d7"),
  1120 => (x"87",x"c7",x"f6",x"c0"),
  1121 => (x"f7",x"f2",x"8e",x"f4"),
  1122 => (x"1e",x"73",x"1e",x"87"),
  1123 => (x"fe",x"49",x"4b",x"71"),
  1124 => (x"49",x"73",x"87",x"c8"),
  1125 => (x"f2",x"87",x"c3",x"fe"),
  1126 => (x"73",x"1e",x"87",x"ea"),
  1127 => (x"c6",x"4b",x"71",x"1e"),
  1128 => (x"c0",x"02",x"4a",x"a3"),
  1129 => (x"8a",x"c1",x"87",x"e3"),
  1130 => (x"8a",x"87",x"d6",x"02"),
  1131 => (x"87",x"e8",x"c1",x"02"),
  1132 => (x"ca",x"c1",x"02",x"8a"),
  1133 => (x"c0",x"02",x"8a",x"87"),
  1134 => (x"02",x"8a",x"87",x"ef"),
  1135 => (x"e9",x"c1",x"87",x"d9"),
  1136 => (x"f6",x"49",x"c7",x"87"),
  1137 => (x"ec",x"c1",x"87",x"c3"),
  1138 => (x"f0",x"da",x"c2",x"87"),
  1139 => (x"c1",x"78",x"df",x"48"),
  1140 => (x"87",x"c1",x"d3",x"49"),
  1141 => (x"c2",x"87",x"de",x"c1"),
  1142 => (x"02",x"bf",x"c8",x"db"),
  1143 => (x"48",x"87",x"cb",x"c1"),
  1144 => (x"db",x"c2",x"88",x"c1"),
  1145 => (x"c1",x"c1",x"58",x"cc"),
  1146 => (x"cc",x"db",x"c2",x"87"),
  1147 => (x"f9",x"c0",x"02",x"bf"),
  1148 => (x"c8",x"db",x"c2",x"87"),
  1149 => (x"80",x"c1",x"48",x"bf"),
  1150 => (x"58",x"cc",x"db",x"c2"),
  1151 => (x"c2",x"87",x"eb",x"c0"),
  1152 => (x"49",x"bf",x"c8",x"db"),
  1153 => (x"db",x"c2",x"89",x"c6"),
  1154 => (x"b7",x"c0",x"59",x"cc"),
  1155 => (x"87",x"da",x"03",x"a9"),
  1156 => (x"48",x"c8",x"db",x"c2"),
  1157 => (x"87",x"d2",x"78",x"c0"),
  1158 => (x"bf",x"cc",x"db",x"c2"),
  1159 => (x"c2",x"87",x"cb",x"02"),
  1160 => (x"48",x"bf",x"c8",x"db"),
  1161 => (x"db",x"c2",x"80",x"c6"),
  1162 => (x"49",x"c0",x"58",x"cc"),
  1163 => (x"73",x"87",x"e6",x"d1"),
  1164 => (x"d6",x"f3",x"c0",x"49"),
  1165 => (x"87",x"cc",x"f0",x"87"),
  1166 => (x"5c",x"5b",x"5e",x"0e"),
  1167 => (x"d4",x"ff",x"0e",x"5d"),
  1168 => (x"59",x"a6",x"dc",x"86"),
  1169 => (x"c0",x"48",x"a6",x"c8"),
  1170 => (x"c1",x"80",x"c4",x"78"),
  1171 => (x"c4",x"78",x"66",x"c0"),
  1172 => (x"c4",x"78",x"c1",x"80"),
  1173 => (x"c2",x"78",x"c1",x"80"),
  1174 => (x"c1",x"48",x"cc",x"db"),
  1175 => (x"f0",x"da",x"c2",x"78"),
  1176 => (x"a8",x"de",x"48",x"bf"),
  1177 => (x"f4",x"87",x"c9",x"05"),
  1178 => (x"a6",x"cc",x"87",x"e6"),
  1179 => (x"87",x"e4",x"cf",x"58"),
  1180 => (x"e4",x"87",x"d0",x"e4"),
  1181 => (x"ff",x"e3",x"87",x"f2"),
  1182 => (x"c0",x"4c",x"70",x"87"),
  1183 => (x"c1",x"02",x"ac",x"fb"),
  1184 => (x"66",x"d8",x"87",x"fb"),
  1185 => (x"87",x"ed",x"c1",x"05"),
  1186 => (x"4a",x"66",x"fc",x"c0"),
  1187 => (x"7e",x"6a",x"82",x"c4"),
  1188 => (x"da",x"c1",x"1e",x"72"),
  1189 => (x"66",x"c4",x"48",x"c9"),
  1190 => (x"4a",x"a1",x"c8",x"49"),
  1191 => (x"aa",x"71",x"41",x"20"),
  1192 => (x"10",x"87",x"f9",x"05"),
  1193 => (x"c0",x"4a",x"26",x"51"),
  1194 => (x"c1",x"48",x"66",x"fc"),
  1195 => (x"6a",x"78",x"d9",x"c3"),
  1196 => (x"74",x"81",x"c7",x"49"),
  1197 => (x"66",x"fc",x"c0",x"51"),
  1198 => (x"c1",x"81",x"c8",x"49"),
  1199 => (x"66",x"fc",x"c0",x"51"),
  1200 => (x"c0",x"81",x"c9",x"49"),
  1201 => (x"66",x"fc",x"c0",x"51"),
  1202 => (x"c0",x"81",x"ca",x"49"),
  1203 => (x"d8",x"1e",x"c1",x"51"),
  1204 => (x"c8",x"49",x"6a",x"1e"),
  1205 => (x"87",x"e4",x"e3",x"81"),
  1206 => (x"c0",x"c1",x"86",x"c8"),
  1207 => (x"a8",x"c0",x"48",x"66"),
  1208 => (x"c8",x"87",x"c7",x"01"),
  1209 => (x"78",x"c1",x"48",x"a6"),
  1210 => (x"c0",x"c1",x"87",x"ce"),
  1211 => (x"88",x"c1",x"48",x"66"),
  1212 => (x"c3",x"58",x"a6",x"d0"),
  1213 => (x"87",x"f0",x"e2",x"87"),
  1214 => (x"c2",x"48",x"a6",x"d0"),
  1215 => (x"02",x"9c",x"74",x"78"),
  1216 => (x"c8",x"87",x"cd",x"cd"),
  1217 => (x"c4",x"c1",x"48",x"66"),
  1218 => (x"cd",x"03",x"a8",x"66"),
  1219 => (x"a6",x"dc",x"87",x"c2"),
  1220 => (x"e8",x"78",x"c0",x"48"),
  1221 => (x"e1",x"78",x"c0",x"80"),
  1222 => (x"4c",x"70",x"87",x"de"),
  1223 => (x"05",x"ac",x"d0",x"c1"),
  1224 => (x"c4",x"87",x"d5",x"c2"),
  1225 => (x"c2",x"e4",x"7e",x"66"),
  1226 => (x"58",x"a6",x"c8",x"87"),
  1227 => (x"70",x"87",x"c9",x"e1"),
  1228 => (x"ac",x"ec",x"c0",x"4c"),
  1229 => (x"87",x"eb",x"c1",x"05"),
  1230 => (x"cb",x"49",x"66",x"c8"),
  1231 => (x"66",x"fc",x"c0",x"91"),
  1232 => (x"4a",x"a1",x"c4",x"81"),
  1233 => (x"a1",x"c8",x"4d",x"6a"),
  1234 => (x"52",x"66",x"c4",x"4a"),
  1235 => (x"79",x"c9",x"fd",x"c0"),
  1236 => (x"70",x"87",x"e5",x"e0"),
  1237 => (x"d8",x"02",x"9c",x"4c"),
  1238 => (x"ac",x"fb",x"c0",x"87"),
  1239 => (x"74",x"87",x"d2",x"02"),
  1240 => (x"87",x"d4",x"e0",x"55"),
  1241 => (x"02",x"9c",x"4c",x"70"),
  1242 => (x"fb",x"c0",x"87",x"c7"),
  1243 => (x"ee",x"ff",x"05",x"ac"),
  1244 => (x"55",x"e0",x"c0",x"87"),
  1245 => (x"c0",x"55",x"c1",x"c2"),
  1246 => (x"66",x"d8",x"7d",x"97"),
  1247 => (x"05",x"a8",x"6e",x"48"),
  1248 => (x"66",x"c8",x"87",x"db"),
  1249 => (x"a8",x"66",x"cc",x"48"),
  1250 => (x"c8",x"87",x"ca",x"04"),
  1251 => (x"80",x"c1",x"48",x"66"),
  1252 => (x"c8",x"58",x"a6",x"cc"),
  1253 => (x"48",x"66",x"cc",x"87"),
  1254 => (x"a6",x"d0",x"88",x"c1"),
  1255 => (x"d7",x"df",x"ff",x"58"),
  1256 => (x"c1",x"4c",x"70",x"87"),
  1257 => (x"c8",x"05",x"ac",x"d0"),
  1258 => (x"48",x"66",x"d4",x"87"),
  1259 => (x"a6",x"d8",x"80",x"c1"),
  1260 => (x"ac",x"d0",x"c1",x"58"),
  1261 => (x"87",x"eb",x"fd",x"02"),
  1262 => (x"d8",x"48",x"66",x"c4"),
  1263 => (x"c9",x"05",x"a8",x"66"),
  1264 => (x"e0",x"c0",x"87",x"e0"),
  1265 => (x"78",x"c0",x"48",x"a6"),
  1266 => (x"fb",x"c0",x"48",x"74"),
  1267 => (x"48",x"7e",x"70",x"88"),
  1268 => (x"e2",x"c9",x"02",x"98"),
  1269 => (x"88",x"cb",x"48",x"87"),
  1270 => (x"98",x"48",x"7e",x"70"),
  1271 => (x"87",x"cd",x"c1",x"02"),
  1272 => (x"70",x"88",x"c9",x"48"),
  1273 => (x"02",x"98",x"48",x"7e"),
  1274 => (x"48",x"87",x"fe",x"c3"),
  1275 => (x"7e",x"70",x"88",x"c4"),
  1276 => (x"ce",x"02",x"98",x"48"),
  1277 => (x"88",x"c1",x"48",x"87"),
  1278 => (x"98",x"48",x"7e",x"70"),
  1279 => (x"87",x"e9",x"c3",x"02"),
  1280 => (x"dc",x"87",x"d6",x"c8"),
  1281 => (x"f0",x"c0",x"48",x"a6"),
  1282 => (x"eb",x"dd",x"ff",x"78"),
  1283 => (x"c0",x"4c",x"70",x"87"),
  1284 => (x"c0",x"02",x"ac",x"ec"),
  1285 => (x"e0",x"c0",x"87",x"c4"),
  1286 => (x"ec",x"c0",x"5c",x"a6"),
  1287 => (x"87",x"cd",x"02",x"ac"),
  1288 => (x"87",x"d4",x"dd",x"ff"),
  1289 => (x"ec",x"c0",x"4c",x"70"),
  1290 => (x"f3",x"ff",x"05",x"ac"),
  1291 => (x"ac",x"ec",x"c0",x"87"),
  1292 => (x"87",x"c4",x"c0",x"02"),
  1293 => (x"87",x"c0",x"dd",x"ff"),
  1294 => (x"1e",x"ca",x"1e",x"c0"),
  1295 => (x"cb",x"49",x"66",x"d0"),
  1296 => (x"66",x"c4",x"c1",x"91"),
  1297 => (x"cc",x"80",x"71",x"48"),
  1298 => (x"66",x"c8",x"58",x"a6"),
  1299 => (x"d0",x"80",x"c4",x"48"),
  1300 => (x"66",x"cc",x"58",x"a6"),
  1301 => (x"dd",x"ff",x"49",x"bf"),
  1302 => (x"1e",x"c1",x"87",x"e2"),
  1303 => (x"66",x"d4",x"1e",x"de"),
  1304 => (x"dd",x"ff",x"49",x"bf"),
  1305 => (x"86",x"d0",x"87",x"d6"),
  1306 => (x"c0",x"48",x"49",x"70"),
  1307 => (x"e8",x"c0",x"88",x"08"),
  1308 => (x"a8",x"c0",x"58",x"a6"),
  1309 => (x"87",x"ee",x"c0",x"06"),
  1310 => (x"48",x"66",x"e4",x"c0"),
  1311 => (x"c0",x"03",x"a8",x"dd"),
  1312 => (x"66",x"c4",x"87",x"e4"),
  1313 => (x"e4",x"c0",x"49",x"bf"),
  1314 => (x"e0",x"c0",x"81",x"66"),
  1315 => (x"66",x"e4",x"c0",x"51"),
  1316 => (x"c4",x"81",x"c1",x"49"),
  1317 => (x"c2",x"81",x"bf",x"66"),
  1318 => (x"e4",x"c0",x"51",x"c1"),
  1319 => (x"81",x"c2",x"49",x"66"),
  1320 => (x"81",x"bf",x"66",x"c4"),
  1321 => (x"48",x"6e",x"51",x"c0"),
  1322 => (x"78",x"d9",x"c3",x"c1"),
  1323 => (x"81",x"c8",x"49",x"6e"),
  1324 => (x"6e",x"51",x"66",x"d0"),
  1325 => (x"d4",x"81",x"c9",x"49"),
  1326 => (x"49",x"6e",x"51",x"66"),
  1327 => (x"66",x"dc",x"81",x"ca"),
  1328 => (x"48",x"66",x"d0",x"51"),
  1329 => (x"a6",x"d4",x"80",x"c1"),
  1330 => (x"48",x"66",x"c8",x"58"),
  1331 => (x"04",x"a8",x"66",x"cc"),
  1332 => (x"c8",x"87",x"cb",x"c0"),
  1333 => (x"80",x"c1",x"48",x"66"),
  1334 => (x"c5",x"58",x"a6",x"cc"),
  1335 => (x"66",x"cc",x"87",x"d9"),
  1336 => (x"d0",x"88",x"c1",x"48"),
  1337 => (x"ce",x"c5",x"58",x"a6"),
  1338 => (x"fe",x"dc",x"ff",x"87"),
  1339 => (x"a6",x"e8",x"c0",x"87"),
  1340 => (x"f6",x"dc",x"ff",x"58"),
  1341 => (x"a6",x"e0",x"c0",x"87"),
  1342 => (x"a8",x"ec",x"c0",x"58"),
  1343 => (x"87",x"ca",x"c0",x"05"),
  1344 => (x"c0",x"48",x"a6",x"dc"),
  1345 => (x"c0",x"78",x"66",x"e4"),
  1346 => (x"d9",x"ff",x"87",x"c4"),
  1347 => (x"66",x"c8",x"87",x"ea"),
  1348 => (x"c0",x"91",x"cb",x"49"),
  1349 => (x"71",x"48",x"66",x"fc"),
  1350 => (x"4a",x"7e",x"70",x"80"),
  1351 => (x"49",x"6e",x"82",x"c8"),
  1352 => (x"e4",x"c0",x"81",x"ca"),
  1353 => (x"66",x"dc",x"51",x"66"),
  1354 => (x"c0",x"81",x"c1",x"49"),
  1355 => (x"c1",x"89",x"66",x"e4"),
  1356 => (x"70",x"30",x"71",x"48"),
  1357 => (x"71",x"89",x"c1",x"49"),
  1358 => (x"de",x"c2",x"7a",x"97"),
  1359 => (x"c0",x"49",x"bf",x"f8"),
  1360 => (x"97",x"29",x"66",x"e4"),
  1361 => (x"71",x"48",x"4a",x"6a"),
  1362 => (x"a6",x"ec",x"c0",x"98"),
  1363 => (x"c4",x"49",x"6e",x"58"),
  1364 => (x"d8",x"4d",x"69",x"81"),
  1365 => (x"66",x"c4",x"48",x"66"),
  1366 => (x"c8",x"c0",x"02",x"a8"),
  1367 => (x"48",x"a6",x"c4",x"87"),
  1368 => (x"c5",x"c0",x"78",x"c0"),
  1369 => (x"48",x"a6",x"c4",x"87"),
  1370 => (x"66",x"c4",x"78",x"c1"),
  1371 => (x"1e",x"e0",x"c0",x"1e"),
  1372 => (x"d9",x"ff",x"49",x"75"),
  1373 => (x"86",x"c8",x"87",x"c6"),
  1374 => (x"b7",x"c0",x"4c",x"70"),
  1375 => (x"d4",x"c1",x"06",x"ac"),
  1376 => (x"c0",x"85",x"74",x"87"),
  1377 => (x"89",x"74",x"49",x"e0"),
  1378 => (x"da",x"c1",x"4b",x"75"),
  1379 => (x"fe",x"71",x"4a",x"d2"),
  1380 => (x"c2",x"87",x"d4",x"ec"),
  1381 => (x"66",x"e0",x"c0",x"85"),
  1382 => (x"c0",x"80",x"c1",x"48"),
  1383 => (x"c0",x"58",x"a6",x"e4"),
  1384 => (x"c1",x"49",x"66",x"e8"),
  1385 => (x"02",x"a9",x"70",x"81"),
  1386 => (x"c4",x"87",x"c8",x"c0"),
  1387 => (x"78",x"c0",x"48",x"a6"),
  1388 => (x"c4",x"87",x"c5",x"c0"),
  1389 => (x"78",x"c1",x"48",x"a6"),
  1390 => (x"c2",x"1e",x"66",x"c4"),
  1391 => (x"e0",x"c0",x"49",x"a4"),
  1392 => (x"70",x"88",x"71",x"48"),
  1393 => (x"49",x"75",x"1e",x"49"),
  1394 => (x"87",x"f0",x"d7",x"ff"),
  1395 => (x"b7",x"c0",x"86",x"c8"),
  1396 => (x"c0",x"ff",x"01",x"a8"),
  1397 => (x"66",x"e0",x"c0",x"87"),
  1398 => (x"87",x"d1",x"c0",x"02"),
  1399 => (x"81",x"c9",x"49",x"6e"),
  1400 => (x"51",x"66",x"e0",x"c0"),
  1401 => (x"c4",x"c1",x"48",x"6e"),
  1402 => (x"cc",x"c0",x"78",x"da"),
  1403 => (x"c9",x"49",x"6e",x"87"),
  1404 => (x"6e",x"51",x"c2",x"81"),
  1405 => (x"c9",x"c6",x"c1",x"48"),
  1406 => (x"48",x"66",x"c8",x"78"),
  1407 => (x"04",x"a8",x"66",x"cc"),
  1408 => (x"c8",x"87",x"cb",x"c0"),
  1409 => (x"80",x"c1",x"48",x"66"),
  1410 => (x"c0",x"58",x"a6",x"cc"),
  1411 => (x"66",x"cc",x"87",x"e9"),
  1412 => (x"d0",x"88",x"c1",x"48"),
  1413 => (x"de",x"c0",x"58",x"a6"),
  1414 => (x"cb",x"d6",x"ff",x"87"),
  1415 => (x"c0",x"4c",x"70",x"87"),
  1416 => (x"c6",x"c1",x"87",x"d5"),
  1417 => (x"c8",x"c0",x"05",x"ac"),
  1418 => (x"48",x"66",x"d0",x"87"),
  1419 => (x"a6",x"d4",x"80",x"c1"),
  1420 => (x"f3",x"d5",x"ff",x"58"),
  1421 => (x"d4",x"4c",x"70",x"87"),
  1422 => (x"80",x"c1",x"48",x"66"),
  1423 => (x"74",x"58",x"a6",x"d8"),
  1424 => (x"cb",x"c0",x"02",x"9c"),
  1425 => (x"48",x"66",x"c8",x"87"),
  1426 => (x"a8",x"66",x"c4",x"c1"),
  1427 => (x"87",x"fe",x"f2",x"04"),
  1428 => (x"87",x"cb",x"d5",x"ff"),
  1429 => (x"c7",x"48",x"66",x"c8"),
  1430 => (x"e5",x"c0",x"03",x"a8"),
  1431 => (x"cc",x"db",x"c2",x"87"),
  1432 => (x"c8",x"78",x"c0",x"48"),
  1433 => (x"91",x"cb",x"49",x"66"),
  1434 => (x"81",x"66",x"fc",x"c0"),
  1435 => (x"6a",x"4a",x"a1",x"c4"),
  1436 => (x"79",x"52",x"c0",x"4a"),
  1437 => (x"c1",x"48",x"66",x"c8"),
  1438 => (x"58",x"a6",x"cc",x"80"),
  1439 => (x"ff",x"04",x"a8",x"c7"),
  1440 => (x"d4",x"ff",x"87",x"db"),
  1441 => (x"f7",x"de",x"ff",x"8e"),
  1442 => (x"61",x"6f",x"4c",x"87"),
  1443 => (x"2e",x"2a",x"20",x"64"),
  1444 => (x"20",x"3a",x"00",x"20"),
  1445 => (x"1e",x"73",x"1e",x"00"),
  1446 => (x"02",x"9b",x"4b",x"71"),
  1447 => (x"db",x"c2",x"87",x"c6"),
  1448 => (x"78",x"c0",x"48",x"c8"),
  1449 => (x"db",x"c2",x"1e",x"c7"),
  1450 => (x"c1",x"1e",x"bf",x"c8"),
  1451 => (x"c2",x"1e",x"fe",x"dd"),
  1452 => (x"49",x"bf",x"f0",x"da"),
  1453 => (x"cc",x"87",x"c1",x"ee"),
  1454 => (x"f0",x"da",x"c2",x"86"),
  1455 => (x"e7",x"e2",x"49",x"bf"),
  1456 => (x"02",x"9b",x"73",x"87"),
  1457 => (x"dd",x"c1",x"87",x"c8"),
  1458 => (x"e2",x"c0",x"49",x"fe"),
  1459 => (x"dd",x"ff",x"87",x"cf"),
  1460 => (x"c1",x"1e",x"87",x"f2"),
  1461 => (x"c0",x"48",x"ea",x"dd"),
  1462 => (x"e1",x"df",x"c1",x"50"),
  1463 => (x"d8",x"ff",x"49",x"bf"),
  1464 => (x"48",x"c0",x"87",x"d2"),
  1465 => (x"c7",x"1e",x"4f",x"26"),
  1466 => (x"49",x"c1",x"87",x"db"),
  1467 => (x"fe",x"87",x"e6",x"fe"),
  1468 => (x"70",x"87",x"f9",x"ee"),
  1469 => (x"87",x"cd",x"02",x"98"),
  1470 => (x"87",x"d3",x"f6",x"fe"),
  1471 => (x"c4",x"02",x"98",x"70"),
  1472 => (x"c2",x"4a",x"c1",x"87"),
  1473 => (x"72",x"4a",x"c0",x"87"),
  1474 => (x"87",x"ce",x"05",x"9a"),
  1475 => (x"dd",x"c1",x"1e",x"c0"),
  1476 => (x"ee",x"c0",x"49",x"c1"),
  1477 => (x"86",x"c4",x"87",x"fa"),
  1478 => (x"db",x"c2",x"87",x"fe"),
  1479 => (x"78",x"c0",x"48",x"c8"),
  1480 => (x"48",x"f0",x"da",x"c2"),
  1481 => (x"c1",x"1e",x"78",x"c0"),
  1482 => (x"c0",x"49",x"cc",x"dd"),
  1483 => (x"c0",x"87",x"e1",x"ee"),
  1484 => (x"87",x"de",x"fe",x"1e"),
  1485 => (x"ee",x"c0",x"49",x"70"),
  1486 => (x"c7",x"c3",x"87",x"d6"),
  1487 => (x"26",x"8e",x"f8",x"87"),
  1488 => (x"20",x"44",x"53",x"4f"),
  1489 => (x"6c",x"69",x"61",x"66"),
  1490 => (x"00",x"2e",x"64",x"65"),
  1491 => (x"74",x"6f",x"6f",x"42"),
  1492 => (x"2e",x"67",x"6e",x"69"),
  1493 => (x"1e",x"00",x"2e",x"2e"),
  1494 => (x"87",x"fe",x"e1",x"c0"),
  1495 => (x"4f",x"26",x"87",x"fa"),
  1496 => (x"87",x"c2",x"fe",x"1e"),
  1497 => (x"48",x"c0",x"87",x"f1"),
  1498 => (x"00",x"00",x"4f",x"26"),
  1499 => (x"00",x"00",x"00",x"01"),
  1500 => (x"78",x"45",x"20",x"80"),
  1501 => (x"80",x"00",x"74",x"69"),
  1502 => (x"63",x"61",x"42",x"20"),
  1503 => (x"0e",x"96",x"00",x"6b"),
  1504 => (x"26",x"dc",x"00",x"00"),
  1505 => (x"00",x"00",x"00",x"00"),
  1506 => (x"00",x"0e",x"96",x"00"),
  1507 => (x"00",x"26",x"fa",x"00"),
  1508 => (x"00",x"00",x"00",x"00"),
  1509 => (x"00",x"00",x"0e",x"96"),
  1510 => (x"00",x"00",x"27",x"18"),
  1511 => (x"96",x"00",x"00",x"00"),
  1512 => (x"36",x"00",x"00",x"0e"),
  1513 => (x"00",x"00",x"00",x"27"),
  1514 => (x"0e",x"96",x"00",x"00"),
  1515 => (x"27",x"54",x"00",x"00"),
  1516 => (x"00",x"00",x"00",x"00"),
  1517 => (x"00",x"0e",x"96",x"00"),
  1518 => (x"00",x"27",x"72",x"00"),
  1519 => (x"00",x"00",x"00",x"00"),
  1520 => (x"00",x"00",x"0e",x"96"),
  1521 => (x"00",x"00",x"27",x"90"),
  1522 => (x"49",x"00",x"00",x"00"),
  1523 => (x"00",x"00",x"00",x"0f"),
  1524 => (x"00",x"00",x"00",x"00"),
  1525 => (x"11",x"9a",x"00",x"00"),
  1526 => (x"00",x"00",x"00",x"00"),
  1527 => (x"00",x"00",x"00",x"00"),
  1528 => (x"00",x"17",x"e5",x"00"),
  1529 => (x"4f",x"4f",x"42",x"00"),
  1530 => (x"20",x"20",x"20",x"54"),
  1531 => (x"4d",x"4f",x"52",x"20"),
  1532 => (x"f0",x"fe",x"1e",x"00"),
  1533 => (x"cd",x"78",x"c0",x"48"),
  1534 => (x"26",x"09",x"79",x"09"),
  1535 => (x"f0",x"fe",x"1e",x"4f"),
  1536 => (x"4f",x"26",x"48",x"bf"),
  1537 => (x"48",x"f0",x"fe",x"1e"),
  1538 => (x"4f",x"26",x"78",x"c1"),
  1539 => (x"48",x"f0",x"fe",x"1e"),
  1540 => (x"4f",x"26",x"78",x"c0"),
  1541 => (x"c0",x"4a",x"71",x"1e"),
  1542 => (x"4f",x"26",x"51",x"52"),
  1543 => (x"5c",x"5b",x"5e",x"0e"),
  1544 => (x"86",x"f4",x"0e",x"5d"),
  1545 => (x"6d",x"97",x"4d",x"71"),
  1546 => (x"4c",x"a5",x"c1",x"7e"),
  1547 => (x"c8",x"48",x"6c",x"97"),
  1548 => (x"48",x"6e",x"58",x"a6"),
  1549 => (x"05",x"a8",x"66",x"c4"),
  1550 => (x"48",x"ff",x"87",x"c5"),
  1551 => (x"ff",x"87",x"e6",x"c0"),
  1552 => (x"a5",x"c2",x"87",x"ca"),
  1553 => (x"4b",x"6c",x"97",x"49"),
  1554 => (x"97",x"4b",x"a3",x"71"),
  1555 => (x"6c",x"97",x"4b",x"6b"),
  1556 => (x"c1",x"48",x"6e",x"7e"),
  1557 => (x"58",x"a6",x"c8",x"80"),
  1558 => (x"a6",x"cc",x"98",x"c7"),
  1559 => (x"7c",x"97",x"70",x"58"),
  1560 => (x"73",x"87",x"e1",x"fe"),
  1561 => (x"26",x"8e",x"f4",x"48"),
  1562 => (x"26",x"4c",x"26",x"4d"),
  1563 => (x"0e",x"4f",x"26",x"4b"),
  1564 => (x"0e",x"5c",x"5b",x"5e"),
  1565 => (x"4c",x"71",x"86",x"f4"),
  1566 => (x"c3",x"4a",x"66",x"d8"),
  1567 => (x"a4",x"c2",x"9a",x"ff"),
  1568 => (x"49",x"6c",x"97",x"4b"),
  1569 => (x"72",x"49",x"a1",x"73"),
  1570 => (x"7e",x"6c",x"97",x"51"),
  1571 => (x"80",x"c1",x"48",x"6e"),
  1572 => (x"c7",x"58",x"a6",x"c8"),
  1573 => (x"58",x"a6",x"cc",x"98"),
  1574 => (x"8e",x"f4",x"54",x"70"),
  1575 => (x"1e",x"87",x"ca",x"ff"),
  1576 => (x"87",x"e8",x"fd",x"1e"),
  1577 => (x"49",x"4a",x"bf",x"e0"),
  1578 => (x"99",x"c0",x"e0",x"c0"),
  1579 => (x"72",x"87",x"cb",x"02"),
  1580 => (x"ee",x"de",x"c2",x"1e"),
  1581 => (x"87",x"f7",x"fe",x"49"),
  1582 => (x"c0",x"fd",x"86",x"c4"),
  1583 => (x"fd",x"7e",x"70",x"87"),
  1584 => (x"26",x"26",x"87",x"c2"),
  1585 => (x"de",x"c2",x"1e",x"4f"),
  1586 => (x"c7",x"fd",x"49",x"ee"),
  1587 => (x"df",x"e2",x"c1",x"87"),
  1588 => (x"87",x"dd",x"fc",x"49"),
  1589 => (x"26",x"87",x"f5",x"c2"),
  1590 => (x"1e",x"73",x"1e",x"4f"),
  1591 => (x"49",x"ee",x"de",x"c2"),
  1592 => (x"70",x"87",x"f9",x"fc"),
  1593 => (x"aa",x"b7",x"c0",x"4a"),
  1594 => (x"87",x"cc",x"c2",x"04"),
  1595 => (x"05",x"aa",x"f0",x"c3"),
  1596 => (x"e6",x"c1",x"87",x"c9"),
  1597 => (x"78",x"c1",x"48",x"c4"),
  1598 => (x"c3",x"87",x"ed",x"c1"),
  1599 => (x"c9",x"05",x"aa",x"e0"),
  1600 => (x"c8",x"e6",x"c1",x"87"),
  1601 => (x"c1",x"78",x"c1",x"48"),
  1602 => (x"e6",x"c1",x"87",x"de"),
  1603 => (x"c6",x"02",x"bf",x"c8"),
  1604 => (x"a2",x"c0",x"c2",x"87"),
  1605 => (x"72",x"87",x"c2",x"4b"),
  1606 => (x"c4",x"e6",x"c1",x"4b"),
  1607 => (x"e0",x"c0",x"02",x"bf"),
  1608 => (x"c4",x"49",x"73",x"87"),
  1609 => (x"c1",x"91",x"29",x"b7"),
  1610 => (x"73",x"81",x"db",x"e7"),
  1611 => (x"c2",x"9a",x"cf",x"4a"),
  1612 => (x"72",x"48",x"c1",x"92"),
  1613 => (x"ff",x"4a",x"70",x"30"),
  1614 => (x"69",x"48",x"72",x"ba"),
  1615 => (x"db",x"79",x"70",x"98"),
  1616 => (x"c4",x"49",x"73",x"87"),
  1617 => (x"c1",x"91",x"29",x"b7"),
  1618 => (x"73",x"81",x"db",x"e7"),
  1619 => (x"c2",x"9a",x"cf",x"4a"),
  1620 => (x"72",x"48",x"c3",x"92"),
  1621 => (x"48",x"4a",x"70",x"30"),
  1622 => (x"79",x"70",x"b0",x"69"),
  1623 => (x"48",x"c8",x"e6",x"c1"),
  1624 => (x"e6",x"c1",x"78",x"c0"),
  1625 => (x"78",x"c0",x"48",x"c4"),
  1626 => (x"49",x"ee",x"de",x"c2"),
  1627 => (x"70",x"87",x"ed",x"fa"),
  1628 => (x"aa",x"b7",x"c0",x"4a"),
  1629 => (x"87",x"f4",x"fd",x"03"),
  1630 => (x"87",x"c4",x"48",x"c0"),
  1631 => (x"4c",x"26",x"4d",x"26"),
  1632 => (x"4f",x"26",x"4b",x"26"),
  1633 => (x"00",x"00",x"00",x"00"),
  1634 => (x"00",x"00",x"00",x"00"),
  1635 => (x"72",x"4a",x"c0",x"1e"),
  1636 => (x"c1",x"91",x"c4",x"49"),
  1637 => (x"c0",x"81",x"db",x"e7"),
  1638 => (x"d0",x"82",x"c1",x"79"),
  1639 => (x"ee",x"04",x"aa",x"b7"),
  1640 => (x"0e",x"4f",x"26",x"87"),
  1641 => (x"5d",x"5c",x"5b",x"5e"),
  1642 => (x"f9",x"4d",x"71",x"0e"),
  1643 => (x"4a",x"75",x"87",x"de"),
  1644 => (x"92",x"2a",x"b7",x"c4"),
  1645 => (x"82",x"db",x"e7",x"c1"),
  1646 => (x"9c",x"cf",x"4c",x"75"),
  1647 => (x"49",x"6a",x"94",x"c2"),
  1648 => (x"c3",x"2b",x"74",x"4b"),
  1649 => (x"74",x"48",x"c2",x"9b"),
  1650 => (x"ff",x"4c",x"70",x"30"),
  1651 => (x"71",x"48",x"74",x"bc"),
  1652 => (x"f8",x"7a",x"70",x"98"),
  1653 => (x"48",x"73",x"87",x"ee"),
  1654 => (x"00",x"87",x"e1",x"fe"),
  1655 => (x"00",x"00",x"00",x"00"),
  1656 => (x"00",x"00",x"00",x"00"),
  1657 => (x"00",x"00",x"00",x"00"),
  1658 => (x"00",x"00",x"00",x"00"),
  1659 => (x"00",x"00",x"00",x"00"),
  1660 => (x"00",x"00",x"00",x"00"),
  1661 => (x"00",x"00",x"00",x"00"),
  1662 => (x"00",x"00",x"00",x"00"),
  1663 => (x"00",x"00",x"00",x"00"),
  1664 => (x"00",x"00",x"00",x"00"),
  1665 => (x"00",x"00",x"00",x"00"),
  1666 => (x"00",x"00",x"00",x"00"),
  1667 => (x"00",x"00",x"00",x"00"),
  1668 => (x"00",x"00",x"00",x"00"),
  1669 => (x"00",x"00",x"00",x"00"),
  1670 => (x"1e",x"00",x"00",x"00"),
  1671 => (x"c8",x"48",x"d0",x"ff"),
  1672 => (x"48",x"71",x"78",x"e1"),
  1673 => (x"78",x"08",x"d4",x"ff"),
  1674 => (x"ff",x"48",x"66",x"c4"),
  1675 => (x"26",x"78",x"08",x"d4"),
  1676 => (x"4a",x"71",x"1e",x"4f"),
  1677 => (x"1e",x"49",x"66",x"c4"),
  1678 => (x"de",x"ff",x"49",x"72"),
  1679 => (x"48",x"d0",x"ff",x"87"),
  1680 => (x"26",x"78",x"e0",x"c0"),
  1681 => (x"73",x"1e",x"4f",x"26"),
  1682 => (x"c8",x"4b",x"71",x"1e"),
  1683 => (x"73",x"1e",x"49",x"66"),
  1684 => (x"a2",x"e0",x"c1",x"4a"),
  1685 => (x"87",x"d9",x"ff",x"49"),
  1686 => (x"26",x"87",x"c4",x"26"),
  1687 => (x"26",x"4c",x"26",x"4d"),
  1688 => (x"1e",x"4f",x"26",x"4b"),
  1689 => (x"4a",x"71",x"1e",x"73"),
  1690 => (x"ab",x"b7",x"c2",x"4b"),
  1691 => (x"a3",x"87",x"c8",x"03"),
  1692 => (x"ff",x"c3",x"4a",x"49"),
  1693 => (x"ce",x"87",x"c7",x"9a"),
  1694 => (x"c3",x"4a",x"49",x"a3"),
  1695 => (x"66",x"c8",x"9a",x"ff"),
  1696 => (x"49",x"72",x"1e",x"49"),
  1697 => (x"26",x"87",x"ea",x"fe"),
  1698 => (x"1e",x"87",x"d4",x"ff"),
  1699 => (x"c3",x"4a",x"d4",x"ff"),
  1700 => (x"d0",x"ff",x"7a",x"ff"),
  1701 => (x"78",x"e1",x"c0",x"48"),
  1702 => (x"de",x"c2",x"7a",x"de"),
  1703 => (x"49",x"7a",x"bf",x"f8"),
  1704 => (x"70",x"28",x"c8",x"48"),
  1705 => (x"d0",x"48",x"71",x"7a"),
  1706 => (x"71",x"7a",x"70",x"28"),
  1707 => (x"70",x"28",x"d8",x"48"),
  1708 => (x"48",x"d0",x"ff",x"7a"),
  1709 => (x"26",x"78",x"e0",x"c0"),
  1710 => (x"d0",x"ff",x"1e",x"4f"),
  1711 => (x"78",x"c9",x"c8",x"48"),
  1712 => (x"d4",x"ff",x"48",x"71"),
  1713 => (x"4f",x"26",x"78",x"08"),
  1714 => (x"49",x"4a",x"71",x"1e"),
  1715 => (x"d0",x"ff",x"87",x"eb"),
  1716 => (x"26",x"78",x"c8",x"48"),
  1717 => (x"1e",x"73",x"1e",x"4f"),
  1718 => (x"df",x"c2",x"4b",x"71"),
  1719 => (x"c3",x"02",x"bf",x"c8"),
  1720 => (x"87",x"eb",x"c2",x"87"),
  1721 => (x"c8",x"48",x"d0",x"ff"),
  1722 => (x"48",x"73",x"78",x"c9"),
  1723 => (x"ff",x"b0",x"e0",x"c0"),
  1724 => (x"c2",x"78",x"08",x"d4"),
  1725 => (x"c0",x"48",x"fc",x"de"),
  1726 => (x"02",x"66",x"c8",x"78"),
  1727 => (x"ff",x"c3",x"87",x"c5"),
  1728 => (x"c0",x"87",x"c2",x"49"),
  1729 => (x"c4",x"df",x"c2",x"49"),
  1730 => (x"02",x"66",x"cc",x"59"),
  1731 => (x"d5",x"c5",x"87",x"c6"),
  1732 => (x"87",x"c4",x"4a",x"d5"),
  1733 => (x"4a",x"ff",x"ff",x"cf"),
  1734 => (x"5a",x"c8",x"df",x"c2"),
  1735 => (x"48",x"c8",x"df",x"c2"),
  1736 => (x"87",x"c4",x"78",x"c1"),
  1737 => (x"4c",x"26",x"4d",x"26"),
  1738 => (x"4f",x"26",x"4b",x"26"),
  1739 => (x"5c",x"5b",x"5e",x"0e"),
  1740 => (x"4a",x"71",x"0e",x"5d"),
  1741 => (x"bf",x"c4",x"df",x"c2"),
  1742 => (x"02",x"9a",x"72",x"4c"),
  1743 => (x"c8",x"49",x"87",x"cb"),
  1744 => (x"cb",x"eb",x"c1",x"91"),
  1745 => (x"c4",x"83",x"71",x"4b"),
  1746 => (x"cb",x"ef",x"c1",x"87"),
  1747 => (x"13",x"4d",x"c0",x"4b"),
  1748 => (x"c2",x"99",x"74",x"49"),
  1749 => (x"48",x"bf",x"c0",x"df"),
  1750 => (x"d4",x"ff",x"b8",x"71"),
  1751 => (x"b7",x"c1",x"78",x"08"),
  1752 => (x"b7",x"c8",x"85",x"2c"),
  1753 => (x"87",x"e7",x"04",x"ad"),
  1754 => (x"bf",x"fc",x"de",x"c2"),
  1755 => (x"c2",x"80",x"c8",x"48"),
  1756 => (x"fe",x"58",x"c0",x"df"),
  1757 => (x"73",x"1e",x"87",x"ee"),
  1758 => (x"13",x"4b",x"71",x"1e"),
  1759 => (x"cb",x"02",x"9a",x"4a"),
  1760 => (x"fe",x"49",x"72",x"87"),
  1761 => (x"4a",x"13",x"87",x"e6"),
  1762 => (x"87",x"f5",x"05",x"9a"),
  1763 => (x"1e",x"87",x"d9",x"fe"),
  1764 => (x"bf",x"fc",x"de",x"c2"),
  1765 => (x"fc",x"de",x"c2",x"49"),
  1766 => (x"78",x"a1",x"c1",x"48"),
  1767 => (x"a9",x"b7",x"c0",x"c4"),
  1768 => (x"ff",x"87",x"db",x"03"),
  1769 => (x"df",x"c2",x"48",x"d4"),
  1770 => (x"c2",x"78",x"bf",x"c0"),
  1771 => (x"49",x"bf",x"fc",x"de"),
  1772 => (x"48",x"fc",x"de",x"c2"),
  1773 => (x"c4",x"78",x"a1",x"c1"),
  1774 => (x"04",x"a9",x"b7",x"c0"),
  1775 => (x"d0",x"ff",x"87",x"e5"),
  1776 => (x"c2",x"78",x"c8",x"48"),
  1777 => (x"c0",x"48",x"c8",x"df"),
  1778 => (x"00",x"4f",x"26",x"78"),
  1779 => (x"00",x"00",x"00",x"00"),
  1780 => (x"00",x"00",x"00",x"00"),
  1781 => (x"5f",x"5f",x"00",x"00"),
  1782 => (x"00",x"00",x"00",x"00"),
  1783 => (x"03",x"00",x"03",x"03"),
  1784 => (x"14",x"00",x"00",x"03"),
  1785 => (x"7f",x"14",x"7f",x"7f"),
  1786 => (x"00",x"00",x"14",x"7f"),
  1787 => (x"6b",x"6b",x"2e",x"24"),
  1788 => (x"4c",x"00",x"12",x"3a"),
  1789 => (x"6c",x"18",x"36",x"6a"),
  1790 => (x"30",x"00",x"32",x"56"),
  1791 => (x"77",x"59",x"4f",x"7e"),
  1792 => (x"00",x"40",x"68",x"3a"),
  1793 => (x"03",x"07",x"04",x"00"),
  1794 => (x"00",x"00",x"00",x"00"),
  1795 => (x"63",x"3e",x"1c",x"00"),
  1796 => (x"00",x"00",x"00",x"41"),
  1797 => (x"3e",x"63",x"41",x"00"),
  1798 => (x"08",x"00",x"00",x"1c"),
  1799 => (x"1c",x"1c",x"3e",x"2a"),
  1800 => (x"00",x"08",x"2a",x"3e"),
  1801 => (x"3e",x"3e",x"08",x"08"),
  1802 => (x"00",x"00",x"08",x"08"),
  1803 => (x"60",x"e0",x"80",x"00"),
  1804 => (x"00",x"00",x"00",x"00"),
  1805 => (x"08",x"08",x"08",x"08"),
  1806 => (x"00",x"00",x"08",x"08"),
  1807 => (x"60",x"60",x"00",x"00"),
  1808 => (x"40",x"00",x"00",x"00"),
  1809 => (x"0c",x"18",x"30",x"60"),
  1810 => (x"00",x"01",x"03",x"06"),
  1811 => (x"4d",x"59",x"7f",x"3e"),
  1812 => (x"00",x"00",x"3e",x"7f"),
  1813 => (x"7f",x"7f",x"06",x"04"),
  1814 => (x"00",x"00",x"00",x"00"),
  1815 => (x"59",x"71",x"63",x"42"),
  1816 => (x"00",x"00",x"46",x"4f"),
  1817 => (x"49",x"49",x"63",x"22"),
  1818 => (x"18",x"00",x"36",x"7f"),
  1819 => (x"7f",x"13",x"16",x"1c"),
  1820 => (x"00",x"00",x"10",x"7f"),
  1821 => (x"45",x"45",x"67",x"27"),
  1822 => (x"00",x"00",x"39",x"7d"),
  1823 => (x"49",x"4b",x"7e",x"3c"),
  1824 => (x"00",x"00",x"30",x"79"),
  1825 => (x"79",x"71",x"01",x"01"),
  1826 => (x"00",x"00",x"07",x"0f"),
  1827 => (x"49",x"49",x"7f",x"36"),
  1828 => (x"00",x"00",x"36",x"7f"),
  1829 => (x"69",x"49",x"4f",x"06"),
  1830 => (x"00",x"00",x"1e",x"3f"),
  1831 => (x"66",x"66",x"00",x"00"),
  1832 => (x"00",x"00",x"00",x"00"),
  1833 => (x"66",x"e6",x"80",x"00"),
  1834 => (x"00",x"00",x"00",x"00"),
  1835 => (x"14",x"14",x"08",x"08"),
  1836 => (x"00",x"00",x"22",x"22"),
  1837 => (x"14",x"14",x"14",x"14"),
  1838 => (x"00",x"00",x"14",x"14"),
  1839 => (x"14",x"14",x"22",x"22"),
  1840 => (x"00",x"00",x"08",x"08"),
  1841 => (x"59",x"51",x"03",x"02"),
  1842 => (x"3e",x"00",x"06",x"0f"),
  1843 => (x"55",x"5d",x"41",x"7f"),
  1844 => (x"00",x"00",x"1e",x"1f"),
  1845 => (x"09",x"09",x"7f",x"7e"),
  1846 => (x"00",x"00",x"7e",x"7f"),
  1847 => (x"49",x"49",x"7f",x"7f"),
  1848 => (x"00",x"00",x"36",x"7f"),
  1849 => (x"41",x"63",x"3e",x"1c"),
  1850 => (x"00",x"00",x"41",x"41"),
  1851 => (x"63",x"41",x"7f",x"7f"),
  1852 => (x"00",x"00",x"1c",x"3e"),
  1853 => (x"49",x"49",x"7f",x"7f"),
  1854 => (x"00",x"00",x"41",x"41"),
  1855 => (x"09",x"09",x"7f",x"7f"),
  1856 => (x"00",x"00",x"01",x"01"),
  1857 => (x"49",x"41",x"7f",x"3e"),
  1858 => (x"00",x"00",x"7a",x"7b"),
  1859 => (x"08",x"08",x"7f",x"7f"),
  1860 => (x"00",x"00",x"7f",x"7f"),
  1861 => (x"7f",x"7f",x"41",x"00"),
  1862 => (x"00",x"00",x"00",x"41"),
  1863 => (x"40",x"40",x"60",x"20"),
  1864 => (x"7f",x"00",x"3f",x"7f"),
  1865 => (x"36",x"1c",x"08",x"7f"),
  1866 => (x"00",x"00",x"41",x"63"),
  1867 => (x"40",x"40",x"7f",x"7f"),
  1868 => (x"7f",x"00",x"40",x"40"),
  1869 => (x"06",x"0c",x"06",x"7f"),
  1870 => (x"7f",x"00",x"7f",x"7f"),
  1871 => (x"18",x"0c",x"06",x"7f"),
  1872 => (x"00",x"00",x"7f",x"7f"),
  1873 => (x"41",x"41",x"7f",x"3e"),
  1874 => (x"00",x"00",x"3e",x"7f"),
  1875 => (x"09",x"09",x"7f",x"7f"),
  1876 => (x"3e",x"00",x"06",x"0f"),
  1877 => (x"7f",x"61",x"41",x"7f"),
  1878 => (x"00",x"00",x"40",x"7e"),
  1879 => (x"19",x"09",x"7f",x"7f"),
  1880 => (x"00",x"00",x"66",x"7f"),
  1881 => (x"59",x"4d",x"6f",x"26"),
  1882 => (x"00",x"00",x"32",x"7b"),
  1883 => (x"7f",x"7f",x"01",x"01"),
  1884 => (x"00",x"00",x"01",x"01"),
  1885 => (x"40",x"40",x"7f",x"3f"),
  1886 => (x"00",x"00",x"3f",x"7f"),
  1887 => (x"70",x"70",x"3f",x"0f"),
  1888 => (x"7f",x"00",x"0f",x"3f"),
  1889 => (x"30",x"18",x"30",x"7f"),
  1890 => (x"41",x"00",x"7f",x"7f"),
  1891 => (x"1c",x"1c",x"36",x"63"),
  1892 => (x"01",x"41",x"63",x"36"),
  1893 => (x"7c",x"7c",x"06",x"03"),
  1894 => (x"61",x"01",x"03",x"06"),
  1895 => (x"47",x"4d",x"59",x"71"),
  1896 => (x"00",x"00",x"41",x"43"),
  1897 => (x"41",x"7f",x"7f",x"00"),
  1898 => (x"01",x"00",x"00",x"41"),
  1899 => (x"18",x"0c",x"06",x"03"),
  1900 => (x"00",x"40",x"60",x"30"),
  1901 => (x"7f",x"41",x"41",x"00"),
  1902 => (x"08",x"00",x"00",x"7f"),
  1903 => (x"06",x"03",x"06",x"0c"),
  1904 => (x"80",x"00",x"08",x"0c"),
  1905 => (x"80",x"80",x"80",x"80"),
  1906 => (x"00",x"00",x"80",x"80"),
  1907 => (x"07",x"03",x"00",x"00"),
  1908 => (x"00",x"00",x"00",x"04"),
  1909 => (x"54",x"54",x"74",x"20"),
  1910 => (x"00",x"00",x"78",x"7c"),
  1911 => (x"44",x"44",x"7f",x"7f"),
  1912 => (x"00",x"00",x"38",x"7c"),
  1913 => (x"44",x"44",x"7c",x"38"),
  1914 => (x"00",x"00",x"00",x"44"),
  1915 => (x"44",x"44",x"7c",x"38"),
  1916 => (x"00",x"00",x"7f",x"7f"),
  1917 => (x"54",x"54",x"7c",x"38"),
  1918 => (x"00",x"00",x"18",x"5c"),
  1919 => (x"05",x"7f",x"7e",x"04"),
  1920 => (x"00",x"00",x"00",x"05"),
  1921 => (x"a4",x"a4",x"bc",x"18"),
  1922 => (x"00",x"00",x"7c",x"fc"),
  1923 => (x"04",x"04",x"7f",x"7f"),
  1924 => (x"00",x"00",x"78",x"7c"),
  1925 => (x"7d",x"3d",x"00",x"00"),
  1926 => (x"00",x"00",x"00",x"40"),
  1927 => (x"fd",x"80",x"80",x"80"),
  1928 => (x"00",x"00",x"00",x"7d"),
  1929 => (x"38",x"10",x"7f",x"7f"),
  1930 => (x"00",x"00",x"44",x"6c"),
  1931 => (x"7f",x"3f",x"00",x"00"),
  1932 => (x"7c",x"00",x"00",x"40"),
  1933 => (x"0c",x"18",x"0c",x"7c"),
  1934 => (x"00",x"00",x"78",x"7c"),
  1935 => (x"04",x"04",x"7c",x"7c"),
  1936 => (x"00",x"00",x"78",x"7c"),
  1937 => (x"44",x"44",x"7c",x"38"),
  1938 => (x"00",x"00",x"38",x"7c"),
  1939 => (x"24",x"24",x"fc",x"fc"),
  1940 => (x"00",x"00",x"18",x"3c"),
  1941 => (x"24",x"24",x"3c",x"18"),
  1942 => (x"00",x"00",x"fc",x"fc"),
  1943 => (x"04",x"04",x"7c",x"7c"),
  1944 => (x"00",x"00",x"08",x"0c"),
  1945 => (x"54",x"54",x"5c",x"48"),
  1946 => (x"00",x"00",x"20",x"74"),
  1947 => (x"44",x"7f",x"3f",x"04"),
  1948 => (x"00",x"00",x"00",x"44"),
  1949 => (x"40",x"40",x"7c",x"3c"),
  1950 => (x"00",x"00",x"7c",x"7c"),
  1951 => (x"60",x"60",x"3c",x"1c"),
  1952 => (x"3c",x"00",x"1c",x"3c"),
  1953 => (x"60",x"30",x"60",x"7c"),
  1954 => (x"44",x"00",x"3c",x"7c"),
  1955 => (x"38",x"10",x"38",x"6c"),
  1956 => (x"00",x"00",x"44",x"6c"),
  1957 => (x"60",x"e0",x"bc",x"1c"),
  1958 => (x"00",x"00",x"1c",x"3c"),
  1959 => (x"5c",x"74",x"64",x"44"),
  1960 => (x"00",x"00",x"44",x"4c"),
  1961 => (x"77",x"3e",x"08",x"08"),
  1962 => (x"00",x"00",x"41",x"41"),
  1963 => (x"7f",x"7f",x"00",x"00"),
  1964 => (x"00",x"00",x"00",x"00"),
  1965 => (x"3e",x"77",x"41",x"41"),
  1966 => (x"02",x"00",x"08",x"08"),
  1967 => (x"02",x"03",x"01",x"01"),
  1968 => (x"7f",x"00",x"01",x"02"),
  1969 => (x"7f",x"7f",x"7f",x"7f"),
  1970 => (x"08",x"00",x"7f",x"7f"),
  1971 => (x"3e",x"1c",x"1c",x"08"),
  1972 => (x"7f",x"7f",x"7f",x"3e"),
  1973 => (x"1c",x"3e",x"3e",x"7f"),
  1974 => (x"00",x"08",x"08",x"1c"),
  1975 => (x"7c",x"7c",x"18",x"10"),
  1976 => (x"00",x"00",x"10",x"18"),
  1977 => (x"7c",x"7c",x"30",x"10"),
  1978 => (x"10",x"00",x"10",x"30"),
  1979 => (x"78",x"60",x"60",x"30"),
  1980 => (x"42",x"00",x"06",x"1e"),
  1981 => (x"3c",x"18",x"3c",x"66"),
  1982 => (x"78",x"00",x"42",x"66"),
  1983 => (x"c6",x"c2",x"6a",x"38"),
  1984 => (x"60",x"00",x"38",x"6c"),
  1985 => (x"00",x"60",x"00",x"00"),
  1986 => (x"0e",x"00",x"60",x"00"),
  1987 => (x"5d",x"5c",x"5b",x"5e"),
  1988 => (x"4c",x"71",x"1e",x"0e"),
  1989 => (x"bf",x"cd",x"df",x"c2"),
  1990 => (x"c0",x"4b",x"c0",x"4d"),
  1991 => (x"02",x"ab",x"74",x"1e"),
  1992 => (x"a6",x"c4",x"87",x"c7"),
  1993 => (x"c5",x"78",x"c0",x"48"),
  1994 => (x"48",x"a6",x"c4",x"87"),
  1995 => (x"66",x"c4",x"78",x"c1"),
  1996 => (x"ee",x"49",x"73",x"1e"),
  1997 => (x"86",x"c8",x"87",x"df"),
  1998 => (x"ef",x"49",x"e0",x"c0"),
  1999 => (x"a5",x"c4",x"87",x"ee"),
  2000 => (x"f0",x"49",x"6a",x"4a"),
  2001 => (x"c6",x"f1",x"87",x"f0"),
  2002 => (x"c1",x"85",x"cb",x"87"),
  2003 => (x"ab",x"b7",x"c8",x"83"),
  2004 => (x"87",x"c7",x"ff",x"04"),
  2005 => (x"26",x"4d",x"26",x"26"),
  2006 => (x"26",x"4b",x"26",x"4c"),
  2007 => (x"4a",x"71",x"1e",x"4f"),
  2008 => (x"5a",x"d1",x"df",x"c2"),
  2009 => (x"48",x"d1",x"df",x"c2"),
  2010 => (x"fe",x"49",x"78",x"c7"),
  2011 => (x"4f",x"26",x"87",x"dd"),
  2012 => (x"71",x"1e",x"73",x"1e"),
  2013 => (x"aa",x"b7",x"c0",x"4a"),
  2014 => (x"c2",x"87",x"d3",x"03"),
  2015 => (x"05",x"bf",x"e9",x"cc"),
  2016 => (x"4b",x"c1",x"87",x"c4"),
  2017 => (x"4b",x"c0",x"87",x"c2"),
  2018 => (x"5b",x"ed",x"cc",x"c2"),
  2019 => (x"cc",x"c2",x"87",x"c4"),
  2020 => (x"cc",x"c2",x"5a",x"ed"),
  2021 => (x"c1",x"4a",x"bf",x"e9"),
  2022 => (x"a2",x"c0",x"c1",x"9a"),
  2023 => (x"87",x"e8",x"ec",x"49"),
  2024 => (x"cc",x"c2",x"48",x"fc"),
  2025 => (x"fe",x"78",x"bf",x"e9"),
  2026 => (x"71",x"1e",x"87",x"ef"),
  2027 => (x"1e",x"66",x"c4",x"4a"),
  2028 => (x"ee",x"ea",x"49",x"72"),
  2029 => (x"4f",x"26",x"26",x"87"),
  2030 => (x"ff",x"4a",x"71",x"1e"),
  2031 => (x"ff",x"c3",x"48",x"d4"),
  2032 => (x"48",x"d0",x"ff",x"78"),
  2033 => (x"ff",x"78",x"e1",x"c0"),
  2034 => (x"78",x"c1",x"48",x"d4"),
  2035 => (x"31",x"c4",x"49",x"72"),
  2036 => (x"d0",x"ff",x"78",x"71"),
  2037 => (x"78",x"e0",x"c0",x"48"),
  2038 => (x"5e",x"0e",x"4f",x"26"),
  2039 => (x"0e",x"5d",x"5c",x"5b"),
  2040 => (x"a6",x"c4",x"86",x"f4"),
  2041 => (x"4b",x"78",x"c0",x"48"),
  2042 => (x"c2",x"7e",x"bf",x"ec"),
  2043 => (x"4d",x"bf",x"cd",x"df"),
  2044 => (x"c2",x"4c",x"bf",x"e8"),
  2045 => (x"49",x"bf",x"e9",x"cc"),
  2046 => (x"cb",x"87",x"de",x"e3"),
  2047 => (x"f0",x"cc",x"49",x"ee"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

