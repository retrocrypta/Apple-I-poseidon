library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"d8dfc287",
    12 => x"86c0c84e",
    13 => x"49d8dfc2",
    14 => x"48d8cdc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087d5dc",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d60299",
    50 => x"c348d4ff",
    51 => x"526878ff",
    52 => x"484966c4",
    53 => x"a6c888c1",
    54 => x"05997158",
    55 => x"4f2687ea",
    56 => x"ff1e731e",
    57 => x"ffc34bd4",
    58 => x"c34a6b7b",
    59 => x"496b7bff",
    60 => x"b17232c8",
    61 => x"6b7bffc3",
    62 => x"7131c84a",
    63 => x"7bffc3b2",
    64 => x"32c8496b",
    65 => x"4871b172",
    66 => x"4d2687c4",
    67 => x"4b264c26",
    68 => x"5e0e4f26",
    69 => x"0e5d5c5b",
    70 => x"d4ff4a71",
    71 => x"c348724c",
    72 => x"7c7098ff",
    73 => x"bfd8cdc2",
    74 => x"d087c805",
    75 => x"30c94866",
    76 => x"d058a6d4",
    77 => x"29d84966",
    78 => x"ffc34871",
    79 => x"d07c7098",
    80 => x"29d04966",
    81 => x"7199ffc3",
    82 => x"4966d07c",
    83 => x"ffc329c8",
    84 => x"d07c7199",
    85 => x"ffc34966",
    86 => x"727c7199",
    87 => x"7129d049",
    88 => x"98ffc348",
    89 => x"4b6c7c70",
    90 => x"4dfff0c9",
    91 => x"05abffc3",
    92 => x"ffc387d0",
    93 => x"c14b6c7c",
    94 => x"87c6028d",
    95 => x"02abffc3",
    96 => x"487387f0",
    97 => x"1e87c3fe",
    98 => x"d4ff49c0",
    99 => x"78ffc348",
   100 => x"c8c381c1",
   101 => x"f104a9b7",
   102 => x"1e4f2687",
   103 => x"87e71e73",
   104 => x"4bdff8c4",
   105 => x"ffc01ec0",
   106 => x"49f7c1f0",
   107 => x"c487e3fd",
   108 => x"05a8c186",
   109 => x"ff87eac0",
   110 => x"ffc348d4",
   111 => x"c0c0c178",
   112 => x"1ec0c0c0",
   113 => x"c1f0e1c0",
   114 => x"c5fd49e9",
   115 => x"7086c487",
   116 => x"87ca0598",
   117 => x"c348d4ff",
   118 => x"48c178ff",
   119 => x"e6fe87cb",
   120 => x"058bc187",
   121 => x"c087fdfe",
   122 => x"87e2fc48",
   123 => x"ff1e731e",
   124 => x"ffc348d4",
   125 => x"c04bd378",
   126 => x"f0ffc01e",
   127 => x"fc49c1c1",
   128 => x"86c487d0",
   129 => x"ca059870",
   130 => x"48d4ff87",
   131 => x"c178ffc3",
   132 => x"fd87cb48",
   133 => x"8bc187f1",
   134 => x"87dbff05",
   135 => x"edfb48c0",
   136 => x"5b5e0e87",
   137 => x"d4ff0e5c",
   138 => x"87dbfd4c",
   139 => x"c01eeac6",
   140 => x"c8c1f0e1",
   141 => x"87dafb49",
   142 => x"a8c186c4",
   143 => x"fe87c802",
   144 => x"48c087ea",
   145 => x"fa87e2c1",
   146 => x"497087d6",
   147 => x"99ffffcf",
   148 => x"02a9eac6",
   149 => x"d3fe87c8",
   150 => x"c148c087",
   151 => x"ffc387cb",
   152 => x"4bf1c07c",
   153 => x"7087f4fc",
   154 => x"ebc00298",
   155 => x"c01ec087",
   156 => x"fac1f0ff",
   157 => x"87dafa49",
   158 => x"987086c4",
   159 => x"c387d905",
   160 => x"496c7cff",
   161 => x"7c7cffc3",
   162 => x"c0c17c7c",
   163 => x"87c40299",
   164 => x"87d548c1",
   165 => x"87d148c0",
   166 => x"c405abc2",
   167 => x"c848c087",
   168 => x"058bc187",
   169 => x"c087fdfe",
   170 => x"87e0f948",
   171 => x"c21e731e",
   172 => x"c148d8cd",
   173 => x"ff4bc778",
   174 => x"78c248d0",
   175 => x"ff87c8fb",
   176 => x"78c348d0",
   177 => x"e5c01ec0",
   178 => x"49c0c1d0",
   179 => x"c487c3f9",
   180 => x"05a8c186",
   181 => x"c24b87c1",
   182 => x"87c505ab",
   183 => x"f9c048c0",
   184 => x"058bc187",
   185 => x"fc87d0ff",
   186 => x"cdc287f7",
   187 => x"987058dc",
   188 => x"c187cd05",
   189 => x"f0ffc01e",
   190 => x"f849d0c1",
   191 => x"86c487d4",
   192 => x"c348d4ff",
   193 => x"fdc278ff",
   194 => x"e0cdc287",
   195 => x"48d0ff58",
   196 => x"d4ff78c2",
   197 => x"78ffc348",
   198 => x"f1f748c1",
   199 => x"5b5e0e87",
   200 => x"710e5d5c",
   201 => x"c54cc04b",
   202 => x"4adfcdee",
   203 => x"c348d4ff",
   204 => x"486878ff",
   205 => x"05a8fec3",
   206 => x"ff87fec0",
   207 => x"9b734dd4",
   208 => x"d087cc02",
   209 => x"49731e66",
   210 => x"c487ecf5",
   211 => x"ff87d686",
   212 => x"d1c448d0",
   213 => x"7dffc378",
   214 => x"c14866d0",
   215 => x"58a6d488",
   216 => x"f0059870",
   217 => x"48d4ff87",
   218 => x"7878ffc3",
   219 => x"c5059b73",
   220 => x"48d0ff87",
   221 => x"4ac178d0",
   222 => x"058ac14c",
   223 => x"7487edfe",
   224 => x"87c6f648",
   225 => x"711e731e",
   226 => x"ff4bc04a",
   227 => x"ffc348d4",
   228 => x"48d0ff78",
   229 => x"ff78c3c4",
   230 => x"ffc348d4",
   231 => x"c01e7278",
   232 => x"d1c1f0ff",
   233 => x"87eaf549",
   234 => x"987086c4",
   235 => x"c887d205",
   236 => x"66cc1ec0",
   237 => x"87e5fd49",
   238 => x"4b7086c4",
   239 => x"c248d0ff",
   240 => x"f5487378",
   241 => x"5e0e87c8",
   242 => x"0e5d5c5b",
   243 => x"ffc01ec0",
   244 => x"49c9c1f0",
   245 => x"d287fbf4",
   246 => x"e0cdc21e",
   247 => x"87fdfc49",
   248 => x"4cc086c8",
   249 => x"b7d284c1",
   250 => x"87f804ac",
   251 => x"97e0cdc2",
   252 => x"c0c349bf",
   253 => x"a9c0c199",
   254 => x"87e7c005",
   255 => x"97e7cdc2",
   256 => x"31d049bf",
   257 => x"97e8cdc2",
   258 => x"32c84abf",
   259 => x"cdc2b172",
   260 => x"4abf97e9",
   261 => x"cf4c71b1",
   262 => x"9cffffff",
   263 => x"34ca84c1",
   264 => x"c287e7c1",
   265 => x"bf97e9cd",
   266 => x"c631c149",
   267 => x"eacdc299",
   268 => x"c74abf97",
   269 => x"b1722ab7",
   270 => x"97e5cdc2",
   271 => x"cf4d4abf",
   272 => x"e6cdc29d",
   273 => x"c34abf97",
   274 => x"c232ca9a",
   275 => x"bf97e7cd",
   276 => x"7333c24b",
   277 => x"e8cdc2b2",
   278 => x"c34bbf97",
   279 => x"b7c69bc0",
   280 => x"c2b2732b",
   281 => x"7148c181",
   282 => x"c1497030",
   283 => x"70307548",
   284 => x"c14c724d",
   285 => x"c8947184",
   286 => x"06adb7c0",
   287 => x"34c187cc",
   288 => x"c0c82db7",
   289 => x"ff01adb7",
   290 => x"487487f4",
   291 => x"0e87fbf1",
   292 => x"5d5c5b5e",
   293 => x"c286f80e",
   294 => x"c048c6d6",
   295 => x"fecdc278",
   296 => x"fb49c01e",
   297 => x"86c487de",
   298 => x"c5059870",
   299 => x"c948c087",
   300 => x"4dc087c0",
   301 => x"edc07ec1",
   302 => x"c249bfe2",
   303 => x"714af4ce",
   304 => x"e4ee4bc8",
   305 => x"05987087",
   306 => x"7ec087c2",
   307 => x"bfdeedc0",
   308 => x"d0cfc249",
   309 => x"4bc8714a",
   310 => x"7087ceee",
   311 => x"87c20598",
   312 => x"026e7ec0",
   313 => x"c287fdc0",
   314 => x"4dbfc4d5",
   315 => x"9ffcd5c2",
   316 => x"c5487ebf",
   317 => x"05a8ead6",
   318 => x"d5c287c7",
   319 => x"ce4dbfc4",
   320 => x"ca486e87",
   321 => x"02a8d5e9",
   322 => x"48c087c5",
   323 => x"c287e3c7",
   324 => x"751efecd",
   325 => x"87ecf949",
   326 => x"987086c4",
   327 => x"c087c505",
   328 => x"87cec748",
   329 => x"bfdeedc0",
   330 => x"d0cfc249",
   331 => x"4bc8714a",
   332 => x"7087f6ec",
   333 => x"87c80598",
   334 => x"48c6d6c2",
   335 => x"87da78c1",
   336 => x"bfe2edc0",
   337 => x"f4cec249",
   338 => x"4bc8714a",
   339 => x"7087daec",
   340 => x"c5c00298",
   341 => x"c648c087",
   342 => x"d5c287d8",
   343 => x"49bf97fc",
   344 => x"05a9d5c1",
   345 => x"c287cdc0",
   346 => x"bf97fdd5",
   347 => x"a9eac249",
   348 => x"87c5c002",
   349 => x"f9c548c0",
   350 => x"fecdc287",
   351 => x"487ebf97",
   352 => x"02a8e9c3",
   353 => x"6e87cec0",
   354 => x"a8ebc348",
   355 => x"87c5c002",
   356 => x"ddc548c0",
   357 => x"c9cec287",
   358 => x"9949bf97",
   359 => x"87ccc005",
   360 => x"97cacec2",
   361 => x"a9c249bf",
   362 => x"87c5c002",
   363 => x"c1c548c0",
   364 => x"cbcec287",
   365 => x"c248bf97",
   366 => x"7058c2d6",
   367 => x"88c1484c",
   368 => x"58c6d6c2",
   369 => x"97cccec2",
   370 => x"817549bf",
   371 => x"97cdcec2",
   372 => x"32c84abf",
   373 => x"c27ea172",
   374 => x"6e48d3da",
   375 => x"cecec278",
   376 => x"c848bf97",
   377 => x"d6c258a6",
   378 => x"c202bfc6",
   379 => x"edc087cf",
   380 => x"c249bfde",
   381 => x"714ad0cf",
   382 => x"ece94bc8",
   383 => x"02987087",
   384 => x"c087c5c0",
   385 => x"87eac348",
   386 => x"bffed5c2",
   387 => x"e7dac24c",
   388 => x"e3cec25c",
   389 => x"c849bf97",
   390 => x"e2cec231",
   391 => x"a14abf97",
   392 => x"e4cec249",
   393 => x"d04abf97",
   394 => x"49a17232",
   395 => x"97e5cec2",
   396 => x"32d84abf",
   397 => x"c449a172",
   398 => x"dac29166",
   399 => x"c281bfd3",
   400 => x"c259dbda",
   401 => x"bf97ebce",
   402 => x"c232c84a",
   403 => x"bf97eace",
   404 => x"c24aa24b",
   405 => x"bf97ecce",
   406 => x"7333d04b",
   407 => x"cec24aa2",
   408 => x"4bbf97ed",
   409 => x"33d89bcf",
   410 => x"c24aa273",
   411 => x"c25adfda",
   412 => x"c292748a",
   413 => x"7248dfda",
   414 => x"c1c178a1",
   415 => x"d0cec287",
   416 => x"c849bf97",
   417 => x"cfcec231",
   418 => x"a14abf97",
   419 => x"c731c549",
   420 => x"29c981ff",
   421 => x"59e7dac2",
   422 => x"97d5cec2",
   423 => x"32c84abf",
   424 => x"97d4cec2",
   425 => x"4aa24bbf",
   426 => x"6e9266c4",
   427 => x"e3dac282",
   428 => x"dbdac25a",
   429 => x"c278c048",
   430 => x"7248d7da",
   431 => x"dac278a1",
   432 => x"dac248e7",
   433 => x"c278bfdb",
   434 => x"c248ebda",
   435 => x"78bfdfda",
   436 => x"bfc6d6c2",
   437 => x"87c9c002",
   438 => x"30c44874",
   439 => x"c9c07e70",
   440 => x"e3dac287",
   441 => x"30c448bf",
   442 => x"d6c27e70",
   443 => x"786e48ca",
   444 => x"8ef848c1",
   445 => x"4c264d26",
   446 => x"4f264b26",
   447 => x"5c5b5e0e",
   448 => x"4a710e5d",
   449 => x"bfc6d6c2",
   450 => x"7287cb02",
   451 => x"722bc74b",
   452 => x"9dffc14d",
   453 => x"4b7287c9",
   454 => x"4d722bc8",
   455 => x"c29dffc3",
   456 => x"83bfd3da",
   457 => x"bfdaedc0",
   458 => x"87d902ab",
   459 => x"5bdeedc0",
   460 => x"1efecdc2",
   461 => x"cbf14973",
   462 => x"7086c487",
   463 => x"87c50598",
   464 => x"e6c048c0",
   465 => x"c6d6c287",
   466 => x"87d202bf",
   467 => x"91c44975",
   468 => x"81fecdc2",
   469 => x"ffcf4c69",
   470 => x"9cffffff",
   471 => x"497587cb",
   472 => x"cdc291c2",
   473 => x"699f81fe",
   474 => x"fe48744c",
   475 => x"5e0e87c6",
   476 => x"0e5d5c5b",
   477 => x"4c7186f8",
   478 => x"87c5059c",
   479 => x"c0c348c0",
   480 => x"7ea4c887",
   481 => x"d878c048",
   482 => x"87c70266",
   483 => x"bf9766d8",
   484 => x"c087c505",
   485 => x"87e9c248",
   486 => x"49c11ec0",
   487 => x"87e3c749",
   488 => x"4d7086c4",
   489 => x"c2c1029d",
   490 => x"ced6c287",
   491 => x"4966d84a",
   492 => x"7087dbe2",
   493 => x"f2c00298",
   494 => x"d84a7587",
   495 => x"4bcb4966",
   496 => x"7087c0e3",
   497 => x"e2c00298",
   498 => x"751ec087",
   499 => x"87c7029d",
   500 => x"c048a6c8",
   501 => x"c887c578",
   502 => x"78c148a6",
   503 => x"c64966c8",
   504 => x"86c487e1",
   505 => x"059d4d70",
   506 => x"7587fefe",
   507 => x"cec1029d",
   508 => x"49a5dc87",
   509 => x"7869486e",
   510 => x"c449a5da",
   511 => x"a4c448a6",
   512 => x"48699f78",
   513 => x"780866c4",
   514 => x"bfc6d6c2",
   515 => x"d487d202",
   516 => x"699f49a5",
   517 => x"ffffc049",
   518 => x"d0487199",
   519 => x"c27e7030",
   520 => x"6e7ec087",
   521 => x"bf66c448",
   522 => x"0866c480",
   523 => x"cc7cc078",
   524 => x"66c449a4",
   525 => x"a4d079bf",
   526 => x"c179c049",
   527 => x"c087c248",
   528 => x"fa8ef848",
   529 => x"5e0e87ee",
   530 => x"710e5c5b",
   531 => x"c1029c4c",
   532 => x"a4c887cb",
   533 => x"c1026949",
   534 => x"496c87c3",
   535 => x"714866cc",
   536 => x"58a6d080",
   537 => x"d6c2b970",
   538 => x"ff4abfc2",
   539 => x"719972ba",
   540 => x"e5c00299",
   541 => x"4ba4c487",
   542 => x"fff9496b",
   543 => x"c27b7087",
   544 => x"49bffed5",
   545 => x"7c71816c",
   546 => x"c2b966cc",
   547 => x"4abfc2d6",
   548 => x"9972baff",
   549 => x"ff059971",
   550 => x"66cc87db",
   551 => x"87d6f97c",
   552 => x"711e731e",
   553 => x"c7029b4b",
   554 => x"49a3c887",
   555 => x"87c50569",
   556 => x"f6c048c0",
   557 => x"d7dac287",
   558 => x"a3c449bf",
   559 => x"c24a6a4a",
   560 => x"fed5c28a",
   561 => x"a17292bf",
   562 => x"c2d6c249",
   563 => x"9a6b4abf",
   564 => x"c049a172",
   565 => x"c859deed",
   566 => x"ea711e66",
   567 => x"86c487e6",
   568 => x"c4059870",
   569 => x"c248c087",
   570 => x"f848c187",
   571 => x"731e87ca",
   572 => x"9b4b711e",
   573 => x"87e4c002",
   574 => x"5bebdac2",
   575 => x"8ac24a73",
   576 => x"bffed5c2",
   577 => x"dac29249",
   578 => x"7248bfd7",
   579 => x"efdac280",
   580 => x"c4487158",
   581 => x"ced6c230",
   582 => x"87edc058",
   583 => x"48e7dac2",
   584 => x"bfdbdac2",
   585 => x"ebdac278",
   586 => x"dfdac248",
   587 => x"d6c278bf",
   588 => x"c902bfc6",
   589 => x"fed5c287",
   590 => x"31c449bf",
   591 => x"dac287c7",
   592 => x"c449bfe3",
   593 => x"ced6c231",
   594 => x"87ecf659",
   595 => x"5c5b5e0e",
   596 => x"c04a710e",
   597 => x"029a724b",
   598 => x"da87e0c0",
   599 => x"699f49a2",
   600 => x"c6d6c24b",
   601 => x"87cf02bf",
   602 => x"9f49a2d4",
   603 => x"c04c4969",
   604 => x"d09cffff",
   605 => x"c087c234",
   606 => x"73b3744c",
   607 => x"87eefd49",
   608 => x"0e87f3f5",
   609 => x"5d5c5b5e",
   610 => x"7186f40e",
   611 => x"727ec04a",
   612 => x"87d8029a",
   613 => x"48facdc2",
   614 => x"cdc278c0",
   615 => x"dac248f2",
   616 => x"c278bfeb",
   617 => x"c248f6cd",
   618 => x"78bfe7da",
   619 => x"48dbd6c2",
   620 => x"d6c250c0",
   621 => x"c249bfca",
   622 => x"4abffacd",
   623 => x"c403aa71",
   624 => x"497287c9",
   625 => x"c00599cf",
   626 => x"edc087e9",
   627 => x"cdc248da",
   628 => x"c278bff2",
   629 => x"c21efecd",
   630 => x"49bff2cd",
   631 => x"48f2cdc2",
   632 => x"7178a1c1",
   633 => x"c487dde6",
   634 => x"d6edc086",
   635 => x"fecdc248",
   636 => x"c087cc78",
   637 => x"48bfd6ed",
   638 => x"c080e0c0",
   639 => x"c258daed",
   640 => x"48bffacd",
   641 => x"cdc280c1",
   642 => x"562758fe",
   643 => x"bf00000b",
   644 => x"9d4dbf97",
   645 => x"87e3c202",
   646 => x"02ade5c3",
   647 => x"c087dcc2",
   648 => x"4bbfd6ed",
   649 => x"1149a3cb",
   650 => x"05accf4c",
   651 => x"7587d2c1",
   652 => x"c199df49",
   653 => x"c291cd89",
   654 => x"c181ced6",
   655 => x"51124aa3",
   656 => x"124aa3c3",
   657 => x"4aa3c551",
   658 => x"a3c75112",
   659 => x"c951124a",
   660 => x"51124aa3",
   661 => x"124aa3ce",
   662 => x"4aa3d051",
   663 => x"a3d25112",
   664 => x"d451124a",
   665 => x"51124aa3",
   666 => x"124aa3d6",
   667 => x"4aa3d851",
   668 => x"a3dc5112",
   669 => x"de51124a",
   670 => x"51124aa3",
   671 => x"fac07ec1",
   672 => x"c8497487",
   673 => x"ebc00599",
   674 => x"d0497487",
   675 => x"87d10599",
   676 => x"c00266dc",
   677 => x"497387cb",
   678 => x"700f66dc",
   679 => x"d3c00298",
   680 => x"c0056e87",
   681 => x"d6c287c6",
   682 => x"50c048ce",
   683 => x"bfd6edc0",
   684 => x"87ddc248",
   685 => x"48dbd6c2",
   686 => x"c27e50c0",
   687 => x"49bfcad6",
   688 => x"bffacdc2",
   689 => x"04aa714a",
   690 => x"c287f7fb",
   691 => x"05bfebda",
   692 => x"c287c8c0",
   693 => x"02bfc6d6",
   694 => x"c287f4c1",
   695 => x"49bff6cd",
   696 => x"c287d9f0",
   697 => x"c458facd",
   698 => x"cdc248a6",
   699 => x"c278bff6",
   700 => x"02bfc6d6",
   701 => x"c487d8c0",
   702 => x"ffcf4966",
   703 => x"99f8ffff",
   704 => x"c5c002a9",
   705 => x"c04cc087",
   706 => x"4cc187e1",
   707 => x"c487dcc0",
   708 => x"ffcf4966",
   709 => x"02a999f8",
   710 => x"c887c8c0",
   711 => x"78c048a6",
   712 => x"c887c5c0",
   713 => x"78c148a6",
   714 => x"744c66c8",
   715 => x"dec0059c",
   716 => x"4966c487",
   717 => x"d5c289c2",
   718 => x"c291bffe",
   719 => x"48bfd7da",
   720 => x"cdc28071",
   721 => x"cdc258f6",
   722 => x"78c048fa",
   723 => x"c087e3f9",
   724 => x"ee8ef448",
   725 => x"000087de",
   726 => x"ffff0000",
   727 => x"0b66ffff",
   728 => x"0b6f0000",
   729 => x"41460000",
   730 => x"20323354",
   731 => x"46002020",
   732 => x"36315441",
   733 => x"00202020",
   734 => x"48d4ff1e",
   735 => x"6878ffc3",
   736 => x"1e4f2648",
   737 => x"c348d4ff",
   738 => x"d0ff78ff",
   739 => x"78e1c048",
   740 => x"d448d4ff",
   741 => x"efdac278",
   742 => x"bfd4ff48",
   743 => x"1e4f2650",
   744 => x"c048d0ff",
   745 => x"4f2678e0",
   746 => x"87ccff1e",
   747 => x"02994970",
   748 => x"fbc087c6",
   749 => x"87f105a9",
   750 => x"4f264871",
   751 => x"5c5b5e0e",
   752 => x"c04b710e",
   753 => x"87f0fe4c",
   754 => x"02994970",
   755 => x"c087f9c0",
   756 => x"c002a9ec",
   757 => x"fbc087f2",
   758 => x"ebc002a9",
   759 => x"b766cc87",
   760 => x"87c703ac",
   761 => x"c20266d0",
   762 => x"71537187",
   763 => x"87c20299",
   764 => x"c3fe84c1",
   765 => x"99497087",
   766 => x"c087cd02",
   767 => x"c702a9ec",
   768 => x"a9fbc087",
   769 => x"87d5ff05",
   770 => x"c30266d0",
   771 => x"7b97c087",
   772 => x"05a9ecc0",
   773 => x"4a7487c4",
   774 => x"4a7487c5",
   775 => x"728a0ac0",
   776 => x"2687c248",
   777 => x"264c264d",
   778 => x"1e4f264b",
   779 => x"7087c9fd",
   780 => x"f0c04a49",
   781 => x"87c904aa",
   782 => x"01aaf9c0",
   783 => x"f0c087c3",
   784 => x"aac1c18a",
   785 => x"c187c904",
   786 => x"c301aada",
   787 => x"8af7c087",
   788 => x"4f264872",
   789 => x"5c5b5e0e",
   790 => x"86f80e5d",
   791 => x"4dc04c71",
   792 => x"c087e0fc",
   793 => x"f3f3c04b",
   794 => x"c049bf97",
   795 => x"87cf04a9",
   796 => x"c187f5fc",
   797 => x"f3f3c083",
   798 => x"ab49bf97",
   799 => x"c087f106",
   800 => x"bf97f3f3",
   801 => x"fb87cf02",
   802 => x"497087ee",
   803 => x"87c60299",
   804 => x"05a9ecc0",
   805 => x"4bc087f1",
   806 => x"7087ddfb",
   807 => x"87d8fb7e",
   808 => x"fb58a6c8",
   809 => x"4a7087d2",
   810 => x"a4c883c1",
   811 => x"49699749",
   812 => x"da05a96e",
   813 => x"49a4c987",
   814 => x"c4496997",
   815 => x"ce05a966",
   816 => x"49a4ca87",
   817 => x"aa496997",
   818 => x"c187c405",
   819 => x"6e87d44d",
   820 => x"a8ecc048",
   821 => x"6e87c802",
   822 => x"a8fbc048",
   823 => x"c087c405",
   824 => x"754dc14b",
   825 => x"effe029d",
   826 => x"87f3fa87",
   827 => x"8ef84873",
   828 => x"0087f0fc",
   829 => x"5c5b5e0e",
   830 => x"86f80e5d",
   831 => x"d4ff7e71",
   832 => x"c21e6e4b",
   833 => x"e949f4da",
   834 => x"86c487e4",
   835 => x"c4029870",
   836 => x"ddc187ea",
   837 => x"6e4dbfec",
   838 => x"87f8fc49",
   839 => x"7058a6c8",
   840 => x"87c50598",
   841 => x"c148a6c4",
   842 => x"48d0ff78",
   843 => x"d5c178c5",
   844 => x"4966c47b",
   845 => x"31c689c1",
   846 => x"97eaddc1",
   847 => x"71484abf",
   848 => x"ff7b70b0",
   849 => x"78c448d0",
   850 => x"97efdac2",
   851 => x"99d049bf",
   852 => x"c587d702",
   853 => x"7bd6c178",
   854 => x"ffc34ac0",
   855 => x"c082c17b",
   856 => x"f504aae0",
   857 => x"48d0ff87",
   858 => x"ffc378c4",
   859 => x"48d0ff7b",
   860 => x"d3c178c5",
   861 => x"c47bc17b",
   862 => x"adb7c078",
   863 => x"87ebc206",
   864 => x"bffcdac2",
   865 => x"029c8d4c",
   866 => x"c287c2c2",
   867 => x"c47efecd",
   868 => x"c0c848a6",
   869 => x"b7c08c78",
   870 => x"87c603ac",
   871 => x"78a4c0c8",
   872 => x"dac24cc0",
   873 => x"49bf97ef",
   874 => x"d00299d0",
   875 => x"c21ec087",
   876 => x"eb49f4da",
   877 => x"86c487ea",
   878 => x"f5c04a70",
   879 => x"fecdc287",
   880 => x"f4dac21e",
   881 => x"87d8eb49",
   882 => x"4a7086c4",
   883 => x"c848d0ff",
   884 => x"d4c178c5",
   885 => x"bf976e7b",
   886 => x"c1486e7b",
   887 => x"c47e7080",
   888 => x"88c14866",
   889 => x"7058a6c8",
   890 => x"e8ff0598",
   891 => x"48d0ff87",
   892 => x"9a7278c4",
   893 => x"c087c505",
   894 => x"87c2c148",
   895 => x"dac21ec1",
   896 => x"c1e949f4",
   897 => x"7486c487",
   898 => x"fefd059c",
   899 => x"adb7c087",
   900 => x"c287d106",
   901 => x"c048f4da",
   902 => x"c080d078",
   903 => x"c280f478",
   904 => x"78bfc0db",
   905 => x"01adb7c0",
   906 => x"ff87d5fd",
   907 => x"78c548d0",
   908 => x"c07bd3c1",
   909 => x"c178c47b",
   910 => x"87c2c048",
   911 => x"8ef848c0",
   912 => x"4c264d26",
   913 => x"4f264b26",
   914 => x"5c5b5e0e",
   915 => x"711e0e5d",
   916 => x"4d4cc04b",
   917 => x"e8c004ab",
   918 => x"d4f1c087",
   919 => x"029d751e",
   920 => x"4ac087c4",
   921 => x"4ac187c2",
   922 => x"d6ec4972",
   923 => x"7086c487",
   924 => x"6e84c17e",
   925 => x"7387c205",
   926 => x"7385c14c",
   927 => x"d8ff06ac",
   928 => x"26486e87",
   929 => x"1e87f9fe",
   930 => x"66c44a71",
   931 => x"7287c505",
   932 => x"87e0f949",
   933 => x"5e0e4f26",
   934 => x"0e5d5c5b",
   935 => x"494c711e",
   936 => x"dbc291de",
   937 => x"85714ddc",
   938 => x"c1026d97",
   939 => x"dbc287dc",
   940 => x"7449bfc8",
   941 => x"cffe7181",
   942 => x"487e7087",
   943 => x"f2c00298",
   944 => x"d0dbc287",
   945 => x"cb4a704b",
   946 => x"dac7ff49",
   947 => x"cb4b7487",
   948 => x"feddc193",
   949 => x"c083c483",
   950 => x"747bcefc",
   951 => x"eac0c149",
   952 => x"c17b7587",
   953 => x"bf97ebdd",
   954 => x"dbc21e49",
   955 => x"d6fe49d0",
   956 => x"7486c487",
   957 => x"d2c0c149",
   958 => x"c149c087",
   959 => x"c287f1c1",
   960 => x"c048f0da",
   961 => x"de49c178",
   962 => x"fc2687cb",
   963 => x"6f4c87f2",
   964 => x"6e696461",
   965 => x"2e2e2e67",
   966 => x"1e731e00",
   967 => x"c2494a71",
   968 => x"81bfc8db",
   969 => x"87e0fc71",
   970 => x"029b4b70",
   971 => x"e84987c4",
   972 => x"dbc287da",
   973 => x"78c048c8",
   974 => x"d8dd49c1",
   975 => x"87c4fc87",
   976 => x"c149c01e",
   977 => x"2687e9c0",
   978 => x"4a711e4f",
   979 => x"c191cb49",
   980 => x"c881fedd",
   981 => x"c2481181",
   982 => x"c258f4da",
   983 => x"c048c8db",
   984 => x"dc49c178",
   985 => x"4f2687ef",
   986 => x"0299711e",
   987 => x"dfc187d2",
   988 => x"50c048d3",
   989 => x"fdc080f7",
   990 => x"ddc140c9",
   991 => x"87ce78f7",
   992 => x"48cfdfc1",
   993 => x"78f0ddc1",
   994 => x"fdc080fc",
   995 => x"4f2678c0",
   996 => x"5c5b5e0e",
   997 => x"86f40e5d",
   998 => x"4dfecdc2",
   999 => x"a6c44cc0",
  1000 => x"c278c048",
  1001 => x"48bfc8db",
  1002 => x"c106a8c0",
  1003 => x"cdc287c0",
  1004 => x"029848fe",
  1005 => x"c087f7c0",
  1006 => x"c81ed4f1",
  1007 => x"87c70266",
  1008 => x"c048a6c4",
  1009 => x"c487c578",
  1010 => x"78c148a6",
  1011 => x"e64966c4",
  1012 => x"86c487f1",
  1013 => x"84c14d70",
  1014 => x"c14866c4",
  1015 => x"58a6c880",
  1016 => x"bfc8dbc2",
  1017 => x"87c603ac",
  1018 => x"ff059d75",
  1019 => x"4cc087c9",
  1020 => x"c3029d75",
  1021 => x"f1c087dc",
  1022 => x"66c81ed4",
  1023 => x"cc87c702",
  1024 => x"78c048a6",
  1025 => x"a6cc87c5",
  1026 => x"cc78c148",
  1027 => x"f2e54966",
  1028 => x"7086c487",
  1029 => x"0298487e",
  1030 => x"4987e4c2",
  1031 => x"699781cb",
  1032 => x"0299d049",
  1033 => x"7487d4c1",
  1034 => x"c191cb49",
  1035 => x"c081fedd",
  1036 => x"c879d9fc",
  1037 => x"51ffc381",
  1038 => x"91de4974",
  1039 => x"4ddcdbc2",
  1040 => x"c1c28571",
  1041 => x"a5c17d97",
  1042 => x"51e0c049",
  1043 => x"97ced6c2",
  1044 => x"87d202bf",
  1045 => x"a5c284c1",
  1046 => x"ced6c24b",
  1047 => x"ff49db4a",
  1048 => x"c187c4c1",
  1049 => x"a5cd87d9",
  1050 => x"c151c049",
  1051 => x"4ba5c284",
  1052 => x"49cb4a6e",
  1053 => x"87efc0ff",
  1054 => x"7487c4c1",
  1055 => x"c191cb49",
  1056 => x"c081fedd",
  1057 => x"c279d6fa",
  1058 => x"bf97ced6",
  1059 => x"7487d802",
  1060 => x"c191de49",
  1061 => x"dcdbc284",
  1062 => x"c283714b",
  1063 => x"dd4aced6",
  1064 => x"c2c0ff49",
  1065 => x"7487d887",
  1066 => x"c293de4b",
  1067 => x"cb83dcdb",
  1068 => x"51c049a3",
  1069 => x"6e7384c1",
  1070 => x"fe49cb4a",
  1071 => x"c487e8ff",
  1072 => x"80c14866",
  1073 => x"c758a6c8",
  1074 => x"c5c003ac",
  1075 => x"fc056e87",
  1076 => x"487487e4",
  1077 => x"e7f58ef4",
  1078 => x"1e731e87",
  1079 => x"cb494b71",
  1080 => x"feddc191",
  1081 => x"4aa1c881",
  1082 => x"48eaddc1",
  1083 => x"a1c95012",
  1084 => x"f3f3c04a",
  1085 => x"ca501248",
  1086 => x"ebddc181",
  1087 => x"c1501148",
  1088 => x"bf97ebdd",
  1089 => x"49c01e49",
  1090 => x"c287fcf5",
  1091 => x"de48f0da",
  1092 => x"d549c178",
  1093 => x"f42687ff",
  1094 => x"5e0e87ea",
  1095 => x"0e5d5c5b",
  1096 => x"4d7186f4",
  1097 => x"c191cb49",
  1098 => x"c881fedd",
  1099 => x"a1ca4aa1",
  1100 => x"48a6c47e",
  1101 => x"bff8dec2",
  1102 => x"bf976e78",
  1103 => x"4866c44b",
  1104 => x"4b702873",
  1105 => x"cc48124c",
  1106 => x"9c7058a6",
  1107 => x"81c984c1",
  1108 => x"b7496997",
  1109 => x"87c204ac",
  1110 => x"976e4cc0",
  1111 => x"66c84abf",
  1112 => x"ff317249",
  1113 => x"9966c4b9",
  1114 => x"30724874",
  1115 => x"71484a70",
  1116 => x"fcdec2b0",
  1117 => x"d2e4c058",
  1118 => x"d449c087",
  1119 => x"497587d7",
  1120 => x"87c7f6c0",
  1121 => x"f7f28ef4",
  1122 => x"1e731e87",
  1123 => x"fe494b71",
  1124 => x"497387c8",
  1125 => x"f287c3fe",
  1126 => x"731e87ea",
  1127 => x"c64b711e",
  1128 => x"c0024aa3",
  1129 => x"8ac187e3",
  1130 => x"8a87d602",
  1131 => x"87e8c102",
  1132 => x"cac1028a",
  1133 => x"c0028a87",
  1134 => x"028a87ef",
  1135 => x"e9c187d9",
  1136 => x"f649c787",
  1137 => x"ecc187c3",
  1138 => x"f0dac287",
  1139 => x"c178df48",
  1140 => x"87c1d349",
  1141 => x"c287dec1",
  1142 => x"02bfc8db",
  1143 => x"4887cbc1",
  1144 => x"dbc288c1",
  1145 => x"c1c158cc",
  1146 => x"ccdbc287",
  1147 => x"f9c002bf",
  1148 => x"c8dbc287",
  1149 => x"80c148bf",
  1150 => x"58ccdbc2",
  1151 => x"c287ebc0",
  1152 => x"49bfc8db",
  1153 => x"dbc289c6",
  1154 => x"b7c059cc",
  1155 => x"87da03a9",
  1156 => x"48c8dbc2",
  1157 => x"87d278c0",
  1158 => x"bfccdbc2",
  1159 => x"c287cb02",
  1160 => x"48bfc8db",
  1161 => x"dbc280c6",
  1162 => x"49c058cc",
  1163 => x"7387e6d1",
  1164 => x"d6f3c049",
  1165 => x"87ccf087",
  1166 => x"5c5b5e0e",
  1167 => x"d4ff0e5d",
  1168 => x"59a6dc86",
  1169 => x"c048a6c8",
  1170 => x"c180c478",
  1171 => x"c47866c0",
  1172 => x"c478c180",
  1173 => x"c278c180",
  1174 => x"c148ccdb",
  1175 => x"f0dac278",
  1176 => x"a8de48bf",
  1177 => x"f487c905",
  1178 => x"a6cc87e6",
  1179 => x"87e4cf58",
  1180 => x"e487d0e4",
  1181 => x"ffe387f2",
  1182 => x"c04c7087",
  1183 => x"c102acfb",
  1184 => x"66d887fb",
  1185 => x"87edc105",
  1186 => x"4a66fcc0",
  1187 => x"7e6a82c4",
  1188 => x"dac11e72",
  1189 => x"66c448c9",
  1190 => x"4aa1c849",
  1191 => x"aa714120",
  1192 => x"1087f905",
  1193 => x"c04a2651",
  1194 => x"c14866fc",
  1195 => x"6a78d9c3",
  1196 => x"7481c749",
  1197 => x"66fcc051",
  1198 => x"c181c849",
  1199 => x"66fcc051",
  1200 => x"c081c949",
  1201 => x"66fcc051",
  1202 => x"c081ca49",
  1203 => x"d81ec151",
  1204 => x"c8496a1e",
  1205 => x"87e4e381",
  1206 => x"c0c186c8",
  1207 => x"a8c04866",
  1208 => x"c887c701",
  1209 => x"78c148a6",
  1210 => x"c0c187ce",
  1211 => x"88c14866",
  1212 => x"c358a6d0",
  1213 => x"87f0e287",
  1214 => x"c248a6d0",
  1215 => x"029c7478",
  1216 => x"c887cdcd",
  1217 => x"c4c14866",
  1218 => x"cd03a866",
  1219 => x"a6dc87c2",
  1220 => x"e878c048",
  1221 => x"e178c080",
  1222 => x"4c7087de",
  1223 => x"05acd0c1",
  1224 => x"c487d5c2",
  1225 => x"c2e47e66",
  1226 => x"58a6c887",
  1227 => x"7087c9e1",
  1228 => x"acecc04c",
  1229 => x"87ebc105",
  1230 => x"cb4966c8",
  1231 => x"66fcc091",
  1232 => x"4aa1c481",
  1233 => x"a1c84d6a",
  1234 => x"5266c44a",
  1235 => x"79c9fdc0",
  1236 => x"7087e5e0",
  1237 => x"d8029c4c",
  1238 => x"acfbc087",
  1239 => x"7487d202",
  1240 => x"87d4e055",
  1241 => x"029c4c70",
  1242 => x"fbc087c7",
  1243 => x"eeff05ac",
  1244 => x"55e0c087",
  1245 => x"c055c1c2",
  1246 => x"66d87d97",
  1247 => x"05a86e48",
  1248 => x"66c887db",
  1249 => x"a866cc48",
  1250 => x"c887ca04",
  1251 => x"80c14866",
  1252 => x"c858a6cc",
  1253 => x"4866cc87",
  1254 => x"a6d088c1",
  1255 => x"d7dfff58",
  1256 => x"c14c7087",
  1257 => x"c805acd0",
  1258 => x"4866d487",
  1259 => x"a6d880c1",
  1260 => x"acd0c158",
  1261 => x"87ebfd02",
  1262 => x"d84866c4",
  1263 => x"c905a866",
  1264 => x"e0c087e0",
  1265 => x"78c048a6",
  1266 => x"fbc04874",
  1267 => x"487e7088",
  1268 => x"e2c90298",
  1269 => x"88cb4887",
  1270 => x"98487e70",
  1271 => x"87cdc102",
  1272 => x"7088c948",
  1273 => x"0298487e",
  1274 => x"4887fec3",
  1275 => x"7e7088c4",
  1276 => x"ce029848",
  1277 => x"88c14887",
  1278 => x"98487e70",
  1279 => x"87e9c302",
  1280 => x"dc87d6c8",
  1281 => x"f0c048a6",
  1282 => x"ebddff78",
  1283 => x"c04c7087",
  1284 => x"c002acec",
  1285 => x"e0c087c4",
  1286 => x"ecc05ca6",
  1287 => x"87cd02ac",
  1288 => x"87d4ddff",
  1289 => x"ecc04c70",
  1290 => x"f3ff05ac",
  1291 => x"acecc087",
  1292 => x"87c4c002",
  1293 => x"87c0ddff",
  1294 => x"1eca1ec0",
  1295 => x"cb4966d0",
  1296 => x"66c4c191",
  1297 => x"cc807148",
  1298 => x"66c858a6",
  1299 => x"d080c448",
  1300 => x"66cc58a6",
  1301 => x"ddff49bf",
  1302 => x"1ec187e2",
  1303 => x"66d41ede",
  1304 => x"ddff49bf",
  1305 => x"86d087d6",
  1306 => x"c0484970",
  1307 => x"e8c08808",
  1308 => x"a8c058a6",
  1309 => x"87eec006",
  1310 => x"4866e4c0",
  1311 => x"c003a8dd",
  1312 => x"66c487e4",
  1313 => x"e4c049bf",
  1314 => x"e0c08166",
  1315 => x"66e4c051",
  1316 => x"c481c149",
  1317 => x"c281bf66",
  1318 => x"e4c051c1",
  1319 => x"81c24966",
  1320 => x"81bf66c4",
  1321 => x"486e51c0",
  1322 => x"78d9c3c1",
  1323 => x"81c8496e",
  1324 => x"6e5166d0",
  1325 => x"d481c949",
  1326 => x"496e5166",
  1327 => x"66dc81ca",
  1328 => x"4866d051",
  1329 => x"a6d480c1",
  1330 => x"4866c858",
  1331 => x"04a866cc",
  1332 => x"c887cbc0",
  1333 => x"80c14866",
  1334 => x"c558a6cc",
  1335 => x"66cc87d9",
  1336 => x"d088c148",
  1337 => x"cec558a6",
  1338 => x"fedcff87",
  1339 => x"a6e8c087",
  1340 => x"f6dcff58",
  1341 => x"a6e0c087",
  1342 => x"a8ecc058",
  1343 => x"87cac005",
  1344 => x"c048a6dc",
  1345 => x"c07866e4",
  1346 => x"d9ff87c4",
  1347 => x"66c887ea",
  1348 => x"c091cb49",
  1349 => x"714866fc",
  1350 => x"4a7e7080",
  1351 => x"496e82c8",
  1352 => x"e4c081ca",
  1353 => x"66dc5166",
  1354 => x"c081c149",
  1355 => x"c18966e4",
  1356 => x"70307148",
  1357 => x"7189c149",
  1358 => x"dec27a97",
  1359 => x"c049bff8",
  1360 => x"972966e4",
  1361 => x"71484a6a",
  1362 => x"a6ecc098",
  1363 => x"c4496e58",
  1364 => x"d84d6981",
  1365 => x"66c44866",
  1366 => x"c8c002a8",
  1367 => x"48a6c487",
  1368 => x"c5c078c0",
  1369 => x"48a6c487",
  1370 => x"66c478c1",
  1371 => x"1ee0c01e",
  1372 => x"d9ff4975",
  1373 => x"86c887c6",
  1374 => x"b7c04c70",
  1375 => x"d4c106ac",
  1376 => x"c0857487",
  1377 => x"897449e0",
  1378 => x"dac14b75",
  1379 => x"fe714ad2",
  1380 => x"c287d4ec",
  1381 => x"66e0c085",
  1382 => x"c080c148",
  1383 => x"c058a6e4",
  1384 => x"c14966e8",
  1385 => x"02a97081",
  1386 => x"c487c8c0",
  1387 => x"78c048a6",
  1388 => x"c487c5c0",
  1389 => x"78c148a6",
  1390 => x"c21e66c4",
  1391 => x"e0c049a4",
  1392 => x"70887148",
  1393 => x"49751e49",
  1394 => x"87f0d7ff",
  1395 => x"b7c086c8",
  1396 => x"c0ff01a8",
  1397 => x"66e0c087",
  1398 => x"87d1c002",
  1399 => x"81c9496e",
  1400 => x"5166e0c0",
  1401 => x"c4c1486e",
  1402 => x"ccc078da",
  1403 => x"c9496e87",
  1404 => x"6e51c281",
  1405 => x"c9c6c148",
  1406 => x"4866c878",
  1407 => x"04a866cc",
  1408 => x"c887cbc0",
  1409 => x"80c14866",
  1410 => x"c058a6cc",
  1411 => x"66cc87e9",
  1412 => x"d088c148",
  1413 => x"dec058a6",
  1414 => x"cbd6ff87",
  1415 => x"c04c7087",
  1416 => x"c6c187d5",
  1417 => x"c8c005ac",
  1418 => x"4866d087",
  1419 => x"a6d480c1",
  1420 => x"f3d5ff58",
  1421 => x"d44c7087",
  1422 => x"80c14866",
  1423 => x"7458a6d8",
  1424 => x"cbc0029c",
  1425 => x"4866c887",
  1426 => x"a866c4c1",
  1427 => x"87fef204",
  1428 => x"87cbd5ff",
  1429 => x"c74866c8",
  1430 => x"e5c003a8",
  1431 => x"ccdbc287",
  1432 => x"c878c048",
  1433 => x"91cb4966",
  1434 => x"8166fcc0",
  1435 => x"6a4aa1c4",
  1436 => x"7952c04a",
  1437 => x"c14866c8",
  1438 => x"58a6cc80",
  1439 => x"ff04a8c7",
  1440 => x"d4ff87db",
  1441 => x"f7deff8e",
  1442 => x"616f4c87",
  1443 => x"2e2a2064",
  1444 => x"203a0020",
  1445 => x"1e731e00",
  1446 => x"029b4b71",
  1447 => x"dbc287c6",
  1448 => x"78c048c8",
  1449 => x"dbc21ec7",
  1450 => x"c11ebfc8",
  1451 => x"c21efedd",
  1452 => x"49bff0da",
  1453 => x"cc87c1ee",
  1454 => x"f0dac286",
  1455 => x"e7e249bf",
  1456 => x"029b7387",
  1457 => x"ddc187c8",
  1458 => x"e2c049fe",
  1459 => x"ddff87cf",
  1460 => x"c11e87f2",
  1461 => x"c048eadd",
  1462 => x"e1dfc150",
  1463 => x"d8ff49bf",
  1464 => x"48c087d2",
  1465 => x"c71e4f26",
  1466 => x"49c187db",
  1467 => x"fe87e6fe",
  1468 => x"7087f9ee",
  1469 => x"87cd0298",
  1470 => x"87d3f6fe",
  1471 => x"c4029870",
  1472 => x"c24ac187",
  1473 => x"724ac087",
  1474 => x"87ce059a",
  1475 => x"ddc11ec0",
  1476 => x"eec049c1",
  1477 => x"86c487fa",
  1478 => x"dbc287fe",
  1479 => x"78c048c8",
  1480 => x"48f0dac2",
  1481 => x"c11e78c0",
  1482 => x"c049ccdd",
  1483 => x"c087e1ee",
  1484 => x"87defe1e",
  1485 => x"eec04970",
  1486 => x"c7c387d6",
  1487 => x"268ef887",
  1488 => x"2044534f",
  1489 => x"6c696166",
  1490 => x"002e6465",
  1491 => x"746f6f42",
  1492 => x"2e676e69",
  1493 => x"1e002e2e",
  1494 => x"87fee1c0",
  1495 => x"4f2687fa",
  1496 => x"87c2fe1e",
  1497 => x"48c087f1",
  1498 => x"00004f26",
  1499 => x"00000001",
  1500 => x"78452080",
  1501 => x"80007469",
  1502 => x"63614220",
  1503 => x"0e96006b",
  1504 => x"26dc0000",
  1505 => x"00000000",
  1506 => x"000e9600",
  1507 => x"0026fa00",
  1508 => x"00000000",
  1509 => x"00000e96",
  1510 => x"00002718",
  1511 => x"96000000",
  1512 => x"3600000e",
  1513 => x"00000027",
  1514 => x"0e960000",
  1515 => x"27540000",
  1516 => x"00000000",
  1517 => x"000e9600",
  1518 => x"00277200",
  1519 => x"00000000",
  1520 => x"00000e96",
  1521 => x"00002790",
  1522 => x"49000000",
  1523 => x"0000000f",
  1524 => x"00000000",
  1525 => x"119a0000",
  1526 => x"00000000",
  1527 => x"00000000",
  1528 => x"0017e500",
  1529 => x"4f4f4200",
  1530 => x"20202054",
  1531 => x"4d4f5220",
  1532 => x"f0fe1e00",
  1533 => x"cd78c048",
  1534 => x"26097909",
  1535 => x"f0fe1e4f",
  1536 => x"4f2648bf",
  1537 => x"48f0fe1e",
  1538 => x"4f2678c1",
  1539 => x"48f0fe1e",
  1540 => x"4f2678c0",
  1541 => x"c04a711e",
  1542 => x"4f265152",
  1543 => x"5c5b5e0e",
  1544 => x"86f40e5d",
  1545 => x"6d974d71",
  1546 => x"4ca5c17e",
  1547 => x"c8486c97",
  1548 => x"486e58a6",
  1549 => x"05a866c4",
  1550 => x"48ff87c5",
  1551 => x"ff87e6c0",
  1552 => x"a5c287ca",
  1553 => x"4b6c9749",
  1554 => x"974ba371",
  1555 => x"6c974b6b",
  1556 => x"c1486e7e",
  1557 => x"58a6c880",
  1558 => x"a6cc98c7",
  1559 => x"7c977058",
  1560 => x"7387e1fe",
  1561 => x"268ef448",
  1562 => x"264c264d",
  1563 => x"0e4f264b",
  1564 => x"0e5c5b5e",
  1565 => x"4c7186f4",
  1566 => x"c34a66d8",
  1567 => x"a4c29aff",
  1568 => x"496c974b",
  1569 => x"7249a173",
  1570 => x"7e6c9751",
  1571 => x"80c1486e",
  1572 => x"c758a6c8",
  1573 => x"58a6cc98",
  1574 => x"8ef45470",
  1575 => x"1e87caff",
  1576 => x"87e8fd1e",
  1577 => x"494abfe0",
  1578 => x"99c0e0c0",
  1579 => x"7287cb02",
  1580 => x"eedec21e",
  1581 => x"87f7fe49",
  1582 => x"c0fd86c4",
  1583 => x"fd7e7087",
  1584 => x"262687c2",
  1585 => x"dec21e4f",
  1586 => x"c7fd49ee",
  1587 => x"dfe2c187",
  1588 => x"87ddfc49",
  1589 => x"2687f5c2",
  1590 => x"1e731e4f",
  1591 => x"49eedec2",
  1592 => x"7087f9fc",
  1593 => x"aab7c04a",
  1594 => x"87ccc204",
  1595 => x"05aaf0c3",
  1596 => x"e6c187c9",
  1597 => x"78c148c4",
  1598 => x"c387edc1",
  1599 => x"c905aae0",
  1600 => x"c8e6c187",
  1601 => x"c178c148",
  1602 => x"e6c187de",
  1603 => x"c602bfc8",
  1604 => x"a2c0c287",
  1605 => x"7287c24b",
  1606 => x"c4e6c14b",
  1607 => x"e0c002bf",
  1608 => x"c4497387",
  1609 => x"c19129b7",
  1610 => x"7381dbe7",
  1611 => x"c29acf4a",
  1612 => x"7248c192",
  1613 => x"ff4a7030",
  1614 => x"694872ba",
  1615 => x"db797098",
  1616 => x"c4497387",
  1617 => x"c19129b7",
  1618 => x"7381dbe7",
  1619 => x"c29acf4a",
  1620 => x"7248c392",
  1621 => x"484a7030",
  1622 => x"7970b069",
  1623 => x"48c8e6c1",
  1624 => x"e6c178c0",
  1625 => x"78c048c4",
  1626 => x"49eedec2",
  1627 => x"7087edfa",
  1628 => x"aab7c04a",
  1629 => x"87f4fd03",
  1630 => x"87c448c0",
  1631 => x"4c264d26",
  1632 => x"4f264b26",
  1633 => x"00000000",
  1634 => x"00000000",
  1635 => x"724ac01e",
  1636 => x"c191c449",
  1637 => x"c081dbe7",
  1638 => x"d082c179",
  1639 => x"ee04aab7",
  1640 => x"0e4f2687",
  1641 => x"5d5c5b5e",
  1642 => x"f94d710e",
  1643 => x"4a7587de",
  1644 => x"922ab7c4",
  1645 => x"82dbe7c1",
  1646 => x"9ccf4c75",
  1647 => x"496a94c2",
  1648 => x"c32b744b",
  1649 => x"7448c29b",
  1650 => x"ff4c7030",
  1651 => x"714874bc",
  1652 => x"f87a7098",
  1653 => x"487387ee",
  1654 => x"0087e1fe",
  1655 => x"00000000",
  1656 => x"00000000",
  1657 => x"00000000",
  1658 => x"00000000",
  1659 => x"00000000",
  1660 => x"00000000",
  1661 => x"00000000",
  1662 => x"00000000",
  1663 => x"00000000",
  1664 => x"00000000",
  1665 => x"00000000",
  1666 => x"00000000",
  1667 => x"00000000",
  1668 => x"00000000",
  1669 => x"00000000",
  1670 => x"1e000000",
  1671 => x"c848d0ff",
  1672 => x"487178e1",
  1673 => x"7808d4ff",
  1674 => x"ff4866c4",
  1675 => x"267808d4",
  1676 => x"4a711e4f",
  1677 => x"1e4966c4",
  1678 => x"deff4972",
  1679 => x"48d0ff87",
  1680 => x"2678e0c0",
  1681 => x"731e4f26",
  1682 => x"c84b711e",
  1683 => x"731e4966",
  1684 => x"a2e0c14a",
  1685 => x"87d9ff49",
  1686 => x"2687c426",
  1687 => x"264c264d",
  1688 => x"1e4f264b",
  1689 => x"4a711e73",
  1690 => x"abb7c24b",
  1691 => x"a387c803",
  1692 => x"ffc34a49",
  1693 => x"ce87c79a",
  1694 => x"c34a49a3",
  1695 => x"66c89aff",
  1696 => x"49721e49",
  1697 => x"2687eafe",
  1698 => x"1e87d4ff",
  1699 => x"c34ad4ff",
  1700 => x"d0ff7aff",
  1701 => x"78e1c048",
  1702 => x"dec27ade",
  1703 => x"497abff8",
  1704 => x"7028c848",
  1705 => x"d048717a",
  1706 => x"717a7028",
  1707 => x"7028d848",
  1708 => x"48d0ff7a",
  1709 => x"2678e0c0",
  1710 => x"d0ff1e4f",
  1711 => x"78c9c848",
  1712 => x"d4ff4871",
  1713 => x"4f267808",
  1714 => x"494a711e",
  1715 => x"d0ff87eb",
  1716 => x"2678c848",
  1717 => x"1e731e4f",
  1718 => x"dfc24b71",
  1719 => x"c302bfc8",
  1720 => x"87ebc287",
  1721 => x"c848d0ff",
  1722 => x"487378c9",
  1723 => x"ffb0e0c0",
  1724 => x"c27808d4",
  1725 => x"c048fcde",
  1726 => x"0266c878",
  1727 => x"ffc387c5",
  1728 => x"c087c249",
  1729 => x"c4dfc249",
  1730 => x"0266cc59",
  1731 => x"d5c587c6",
  1732 => x"87c44ad5",
  1733 => x"4affffcf",
  1734 => x"5ac8dfc2",
  1735 => x"48c8dfc2",
  1736 => x"87c478c1",
  1737 => x"4c264d26",
  1738 => x"4f264b26",
  1739 => x"5c5b5e0e",
  1740 => x"4a710e5d",
  1741 => x"bfc4dfc2",
  1742 => x"029a724c",
  1743 => x"c84987cb",
  1744 => x"cbebc191",
  1745 => x"c483714b",
  1746 => x"cbefc187",
  1747 => x"134dc04b",
  1748 => x"c2997449",
  1749 => x"48bfc0df",
  1750 => x"d4ffb871",
  1751 => x"b7c17808",
  1752 => x"b7c8852c",
  1753 => x"87e704ad",
  1754 => x"bffcdec2",
  1755 => x"c280c848",
  1756 => x"fe58c0df",
  1757 => x"731e87ee",
  1758 => x"134b711e",
  1759 => x"cb029a4a",
  1760 => x"fe497287",
  1761 => x"4a1387e6",
  1762 => x"87f5059a",
  1763 => x"1e87d9fe",
  1764 => x"bffcdec2",
  1765 => x"fcdec249",
  1766 => x"78a1c148",
  1767 => x"a9b7c0c4",
  1768 => x"ff87db03",
  1769 => x"dfc248d4",
  1770 => x"c278bfc0",
  1771 => x"49bffcde",
  1772 => x"48fcdec2",
  1773 => x"c478a1c1",
  1774 => x"04a9b7c0",
  1775 => x"d0ff87e5",
  1776 => x"c278c848",
  1777 => x"c048c8df",
  1778 => x"004f2678",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"5f5f0000",
  1782 => x"00000000",
  1783 => x"03000303",
  1784 => x"14000003",
  1785 => x"7f147f7f",
  1786 => x"0000147f",
  1787 => x"6b6b2e24",
  1788 => x"4c00123a",
  1789 => x"6c18366a",
  1790 => x"30003256",
  1791 => x"77594f7e",
  1792 => x"0040683a",
  1793 => x"03070400",
  1794 => x"00000000",
  1795 => x"633e1c00",
  1796 => x"00000041",
  1797 => x"3e634100",
  1798 => x"0800001c",
  1799 => x"1c1c3e2a",
  1800 => x"00082a3e",
  1801 => x"3e3e0808",
  1802 => x"00000808",
  1803 => x"60e08000",
  1804 => x"00000000",
  1805 => x"08080808",
  1806 => x"00000808",
  1807 => x"60600000",
  1808 => x"40000000",
  1809 => x"0c183060",
  1810 => x"00010306",
  1811 => x"4d597f3e",
  1812 => x"00003e7f",
  1813 => x"7f7f0604",
  1814 => x"00000000",
  1815 => x"59716342",
  1816 => x"0000464f",
  1817 => x"49496322",
  1818 => x"1800367f",
  1819 => x"7f13161c",
  1820 => x"0000107f",
  1821 => x"45456727",
  1822 => x"0000397d",
  1823 => x"494b7e3c",
  1824 => x"00003079",
  1825 => x"79710101",
  1826 => x"0000070f",
  1827 => x"49497f36",
  1828 => x"0000367f",
  1829 => x"69494f06",
  1830 => x"00001e3f",
  1831 => x"66660000",
  1832 => x"00000000",
  1833 => x"66e68000",
  1834 => x"00000000",
  1835 => x"14140808",
  1836 => x"00002222",
  1837 => x"14141414",
  1838 => x"00001414",
  1839 => x"14142222",
  1840 => x"00000808",
  1841 => x"59510302",
  1842 => x"3e00060f",
  1843 => x"555d417f",
  1844 => x"00001e1f",
  1845 => x"09097f7e",
  1846 => x"00007e7f",
  1847 => x"49497f7f",
  1848 => x"0000367f",
  1849 => x"41633e1c",
  1850 => x"00004141",
  1851 => x"63417f7f",
  1852 => x"00001c3e",
  1853 => x"49497f7f",
  1854 => x"00004141",
  1855 => x"09097f7f",
  1856 => x"00000101",
  1857 => x"49417f3e",
  1858 => x"00007a7b",
  1859 => x"08087f7f",
  1860 => x"00007f7f",
  1861 => x"7f7f4100",
  1862 => x"00000041",
  1863 => x"40406020",
  1864 => x"7f003f7f",
  1865 => x"361c087f",
  1866 => x"00004163",
  1867 => x"40407f7f",
  1868 => x"7f004040",
  1869 => x"060c067f",
  1870 => x"7f007f7f",
  1871 => x"180c067f",
  1872 => x"00007f7f",
  1873 => x"41417f3e",
  1874 => x"00003e7f",
  1875 => x"09097f7f",
  1876 => x"3e00060f",
  1877 => x"7f61417f",
  1878 => x"0000407e",
  1879 => x"19097f7f",
  1880 => x"0000667f",
  1881 => x"594d6f26",
  1882 => x"0000327b",
  1883 => x"7f7f0101",
  1884 => x"00000101",
  1885 => x"40407f3f",
  1886 => x"00003f7f",
  1887 => x"70703f0f",
  1888 => x"7f000f3f",
  1889 => x"3018307f",
  1890 => x"41007f7f",
  1891 => x"1c1c3663",
  1892 => x"01416336",
  1893 => x"7c7c0603",
  1894 => x"61010306",
  1895 => x"474d5971",
  1896 => x"00004143",
  1897 => x"417f7f00",
  1898 => x"01000041",
  1899 => x"180c0603",
  1900 => x"00406030",
  1901 => x"7f414100",
  1902 => x"0800007f",
  1903 => x"0603060c",
  1904 => x"8000080c",
  1905 => x"80808080",
  1906 => x"00008080",
  1907 => x"07030000",
  1908 => x"00000004",
  1909 => x"54547420",
  1910 => x"0000787c",
  1911 => x"44447f7f",
  1912 => x"0000387c",
  1913 => x"44447c38",
  1914 => x"00000044",
  1915 => x"44447c38",
  1916 => x"00007f7f",
  1917 => x"54547c38",
  1918 => x"0000185c",
  1919 => x"057f7e04",
  1920 => x"00000005",
  1921 => x"a4a4bc18",
  1922 => x"00007cfc",
  1923 => x"04047f7f",
  1924 => x"0000787c",
  1925 => x"7d3d0000",
  1926 => x"00000040",
  1927 => x"fd808080",
  1928 => x"0000007d",
  1929 => x"38107f7f",
  1930 => x"0000446c",
  1931 => x"7f3f0000",
  1932 => x"7c000040",
  1933 => x"0c180c7c",
  1934 => x"0000787c",
  1935 => x"04047c7c",
  1936 => x"0000787c",
  1937 => x"44447c38",
  1938 => x"0000387c",
  1939 => x"2424fcfc",
  1940 => x"0000183c",
  1941 => x"24243c18",
  1942 => x"0000fcfc",
  1943 => x"04047c7c",
  1944 => x"0000080c",
  1945 => x"54545c48",
  1946 => x"00002074",
  1947 => x"447f3f04",
  1948 => x"00000044",
  1949 => x"40407c3c",
  1950 => x"00007c7c",
  1951 => x"60603c1c",
  1952 => x"3c001c3c",
  1953 => x"6030607c",
  1954 => x"44003c7c",
  1955 => x"3810386c",
  1956 => x"0000446c",
  1957 => x"60e0bc1c",
  1958 => x"00001c3c",
  1959 => x"5c746444",
  1960 => x"0000444c",
  1961 => x"773e0808",
  1962 => x"00004141",
  1963 => x"7f7f0000",
  1964 => x"00000000",
  1965 => x"3e774141",
  1966 => x"02000808",
  1967 => x"02030101",
  1968 => x"7f000102",
  1969 => x"7f7f7f7f",
  1970 => x"08007f7f",
  1971 => x"3e1c1c08",
  1972 => x"7f7f7f3e",
  1973 => x"1c3e3e7f",
  1974 => x"0008081c",
  1975 => x"7c7c1810",
  1976 => x"00001018",
  1977 => x"7c7c3010",
  1978 => x"10001030",
  1979 => x"78606030",
  1980 => x"4200061e",
  1981 => x"3c183c66",
  1982 => x"78004266",
  1983 => x"c6c26a38",
  1984 => x"6000386c",
  1985 => x"00600000",
  1986 => x"0e006000",
  1987 => x"5d5c5b5e",
  1988 => x"4c711e0e",
  1989 => x"bfcddfc2",
  1990 => x"c04bc04d",
  1991 => x"02ab741e",
  1992 => x"a6c487c7",
  1993 => x"c578c048",
  1994 => x"48a6c487",
  1995 => x"66c478c1",
  1996 => x"ee49731e",
  1997 => x"86c887df",
  1998 => x"ef49e0c0",
  1999 => x"a5c487ee",
  2000 => x"f0496a4a",
  2001 => x"c6f187f0",
  2002 => x"c185cb87",
  2003 => x"abb7c883",
  2004 => x"87c7ff04",
  2005 => x"264d2626",
  2006 => x"264b264c",
  2007 => x"4a711e4f",
  2008 => x"5ad1dfc2",
  2009 => x"48d1dfc2",
  2010 => x"fe4978c7",
  2011 => x"4f2687dd",
  2012 => x"711e731e",
  2013 => x"aab7c04a",
  2014 => x"c287d303",
  2015 => x"05bfe9cc",
  2016 => x"4bc187c4",
  2017 => x"4bc087c2",
  2018 => x"5bedccc2",
  2019 => x"ccc287c4",
  2020 => x"ccc25aed",
  2021 => x"c14abfe9",
  2022 => x"a2c0c19a",
  2023 => x"87e8ec49",
  2024 => x"ccc248fc",
  2025 => x"fe78bfe9",
  2026 => x"711e87ef",
  2027 => x"1e66c44a",
  2028 => x"eeea4972",
  2029 => x"4f262687",
  2030 => x"ff4a711e",
  2031 => x"ffc348d4",
  2032 => x"48d0ff78",
  2033 => x"ff78e1c0",
  2034 => x"78c148d4",
  2035 => x"31c44972",
  2036 => x"d0ff7871",
  2037 => x"78e0c048",
  2038 => x"5e0e4f26",
  2039 => x"0e5d5c5b",
  2040 => x"a6c486f4",
  2041 => x"4b78c048",
  2042 => x"c27ebfec",
  2043 => x"4dbfcddf",
  2044 => x"c24cbfe8",
  2045 => x"49bfe9cc",
  2046 => x"cb87dee3",
  2047 => x"f0cc49ee",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
